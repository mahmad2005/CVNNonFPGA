library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


package nn_package is

    -- Network architecture parameters
    constant NUM_X : integer := 128; -- Number of inputs
    constant NUM_L1 : integer := 20; -- Number of hidden layer neurons
    constant NUM_Y : integer := 10; -- Number of outputs
    
    constant BATCH_SIZE : integer := 16; -- Input batch size
    constant NUMBER_OF_BATCH : integer := 8; --Number of batch 

    -- Data representation constants
    constant N : integer := 16; -- Number of bits (data width) 32
    constant F : integer := 8; -- Number of fractional bits 20
    constant I : integer := N-F; -- Number of integer bits
    constant ONE : real := 2.0**F;
    constant ONE_int : integer := integer(ONE); -- 1 in fixed point representation

    -- Array types (for representing signals throughout the network
    type x_array is array(0 to NUM_X-1) of signed(N-1 downto 0); -- Array of inputs
    type y_array is array(0 to NUM_Y-1) of signed(N-1 downto 0); -- Array of outputs
    type sum1_array is array(0 to NUM_L1-1) of signed(N-1 downto 0); -- Array of hidden neuron outputs
    type sum2_array is array(0 to NUM_Y-1) of signed(N-1 downto 0); -- Array of output neuron outputs
    type a_array is array(0 to NUM_L1-1) of signed(N-1 downto 0); -- Array of hidden activation function outputs
    
    type batch_x_array is array(0 to BATCH_SIZE-1) of signed(N-1 downto 0); -- Array of input_batch

    -- Array types (real valued for representation of bias, weight and
    -- normalization parameters
    type b1r_array is array(0 to NUM_L1-1) of real; -- Hidden layer biases
    type b2r_array is array(0 to NUM_Y-1) of real; -- Output layer biases
    type w1r_array is array(0 to NUM_X*NUM_L1-1) of real; -- Hidden layer weights
    type w2r_array is array(0 to NUM_L1*NUM_Y-1) of real; -- Output layer weights
    type p1r_array is array(0 to NUM_X-1) of real; -- Normalization parameters
    type p2r_array is array(0 to NUM_Y-1) of real; -- Denormalization parameters

    -- Array types (signed valued for representation of bias, weight and
    -- normalization parameters
    type b1_array is array (0 to NUM_L1-1) of signed(N-1 downto 0); -- Hidden layer biases
    type b2_array is array (0 to NUM_Y-1) of signed(N-1 downto 0); -- Output layer biases
    type w1_array is array (0 to NUM_L1-1) of x_array; -- Hidden layer weights
    type w2_array is array (0 to NUM_Y-1) of a_array; -- Output layer weights
    type p1_array is array (0 to NUM_X-1) of signed(N-1 downto 0); -- Normalization parameters
    type p2_array is array (0 to NUM_Y-1) of signed(N-1 downto 0); -- Denormalization parameters

    type input_array is array(0 to 127) of real;-- input array
    type output_array is array(0 to 127) of real;-- output array
    -- Real weights and biases
    -- hidden layer biases
    constant b1r : b1r_array := (-1.035337448120117188e+01,-1.897765040397644043e+00,-1.920840859413146973e+00,-2.359372854232788086e+00,-1.115016460418701172e+00,-1.088147163391113281e+00,2.012675285339355469e+00,-2.423217058181762695e+00,-6.122645378112792969e+00,1.245750069618225098e+00,-1.218131542205810547e+01,-1.310552358627319336e-01,7.056146860122680664e-01,2.195918560028076172e+00,-1.561551856994628906e+01,-5.849385857582092285e-01,-1.243088483810424805e+00,-1.523425674438476562e+01,3.293507337570190430e+00,1.068536520004272461e+00);
    constant b1r_imag : b1r_array := (-1.921094894409179688e+00,-1.460755443572998047e+01,-1.007697677612304688e+01,-1.070056247711181641e+01,-8.666425704956054688e+00,-3.615695238113403320e+00,-1.000465679168701172e+01,-7.189449310302734375e+00,-4.318104386329650879e-01,-1.181687927246093750e+01,1.109672665596008301e+00,-1.826949501037597656e+01,-1.105520820617675781e+01,-9.796757698059082031e+00,9.170024394989013672e-01,-1.672972869873046875e+01,-8.574002265930175781e+00,1.287263035774230957e+00,-5.433824062347412109e+00,-1.365888309478759766e+01);
    constant b2r : b2r_array := (-2.067325353622436523e+00,3.398120105266571045e-01,1.806251287460327148e+00,-1.384781241416931152e+00,9.496596455574035645e-01,-7.700572609901428223e-01,-6.157314777374267578e-01,1.061525382101535797e-02,-3.295247554779052734e-01,2.132420301437377930e+00);
    constant b2r_imag : b2r_array := (-2.150891542434692383e+00,7.976756691932678223e-01,1.943687438964843750e+00,-1.297501802444458008e+00,9.918466806411743164e-01,-9.170073866844177246e-01,-1.103455543518066406e+00,-2.379931360483169556e-01,-3.311586081981658936e-01,2.218790292739868164e+00);
    -- hidden layer weights
    constant w1r : w1r_array := (-3.901882171630859375e-01,4.011066630482673645e-02,2.853605151176452637e-01,2.956728450953960419e-02,-2.371521890163421631e-01,3.665456771850585938e-01,2.379177361726760864e-01,1.301534622907638550e-01,5.603278279304504395e-01,5.642318129539489746e-01,3.316210582852363586e-02,-1.418123990297317505e-01,4.084816277027130127e-01,2.449025660753250122e-01,9.050515480339527130e-03,2.381803542375564575e-01,3.286333084106445312e-01,1.010095402598381042e-01,2.018356323242187500e-01,1.469336152076721191e-01,-4.135400429368019104e-02,1.406012475490570068e-01,4.228760004043579102e-01,-3.554078564047813416e-02,-2.499116212129592896e-02,2.184367328882217407e-01,5.037612840533256531e-02,3.428683578968048096e-01,-1.676139235496520996e-01,4.672779142856597900e-02,1.974488943815231323e-01,-7.830626517534255981e-02,-1.466420441865921021e-01,1.512339562177658081e-01,-6.111425906419754028e-02,9.858278930187225342e-02,-3.922166768461465836e-03,2.226373851299285889e-01,2.221276462078094482e-01,-2.926456928253173828e-02,1.489930506795644760e-02,2.286541908979415894e-01,-8.930214494466781616e-02,1.942093372344970703e-01,3.465779125690460205e-01,6.171369552612304688e-02,1.639578044414520264e-01,-4.247864708304405212e-02,1.658212989568710327e-01,3.038277849555015564e-02,1.004301607608795166e-01,-2.915490977466106415e-02,5.906284227967262268e-02,1.029444113373756409e-01,-2.756047435104846954e-02,2.621888816356658936e-01,-7.680781930685043335e-02,-5.357276275753974915e-02,1.876520216464996338e-01,1.332043949514627457e-02,3.090025782585144043e-01,-1.260142177343368530e-01,-8.009829372167587280e-02,-1.310102939605712891e-01,2.438536100089550018e-02,6.549530476331710815e-02,4.735121503472328186e-02,4.972156137228012085e-02,-4.392556473612785339e-02,-8.166747540235519409e-02,-1.396718472242355347e-01,1.041515767574310303e-01,-3.446754813194274902e-02,-1.196118742227554321e-01,1.746238023042678833e-02,1.867916733026504517e-01,1.207171380519866943e-01,-1.301623582839965820e-01,-1.208146214485168457e-01,-5.879015102982521057e-02,5.855090543627738953e-02,-2.937852442264556885e-01,-3.708827309310436249e-03,-3.196318149566650391e-01,-2.419763803482055664e-02,-6.870904564857482910e-02,6.651479005813598633e-02,3.379221260547637939e-01,-1.305372565984725952e-01,-3.360483795404434204e-02,1.502999812364578247e-01,-1.541787832975387573e-01,-9.780462831258773804e-02,-1.958019137382507324e-01,-1.091033816337585449e-01,1.753643341362476349e-02,-7.492101937532424927e-02,7.486672699451446533e-02,-9.826976805925369263e-02,-1.658490002155303955e-01,2.313251346349716187e-01,6.108615081757307053e-03,-9.776693582534790039e-02,9.378809481859207153e-02,-1.434611678123474121e-01,1.682232022285461426e-01,-4.302910342812538147e-02,-1.184836179018020630e-01,1.989995688199996948e-02,3.912518322467803955e-01,-1.782655417919158936e-01,-7.291361689567565918e-02,3.514314889907836914e-01,1.098189800977706909e-01,1.223654523491859436e-01,4.594437479972839355e-01,1.225606575608253479e-01,-6.065908446907997131e-02,1.702614873647689819e-01,2.713257372379302979e-01,-2.419094294309616089e-01,-2.055377513170242310e-01,-2.389217764139175415e-01,-1.080402582883834839e-01,6.975372135639190674e-02,1.849393360316753387e-02,4.812907576560974121e-01,4.251812398433685303e-02,-3.485269546508789062e-01,-2.892071604728698730e-01,-1.793103516101837158e-01,-1.168701946735382080e-01,-5.659558176994323730e-01,-1.607301086187362671e-01,2.206217497587203979e-01,2.389220297336578369e-01,2.321081757545471191e-01,1.909483373165130615e-01,3.794648125767707825e-02,-3.755543380975723267e-02,-4.885422997176647186e-03,5.741427466273307800e-02,1.076057404279708862e-01,9.243579208850860596e-02,1.240135952830314636e-01,3.924762830138206482e-02,2.340009957551956177e-01,-1.122059747576713562e-01,-8.787113474681973457e-04,5.953956767916679382e-02,-5.528088659048080444e-02,2.018535733222961426e-01,1.071153134107589722e-01,3.414735943078994751e-02,1.442320942878723145e-01,1.963927000761032104e-01,6.819085776805877686e-02,2.765402197837829590e-01,1.270516365766525269e-01,1.700378209352493286e-01,8.131939917802810669e-02,8.897923678159713745e-02,7.168569415807723999e-02,5.550422891974449158e-02,1.627590060234069824e-01,1.489408314228057861e-01,1.226608604192733765e-01,5.173910036683082581e-02,1.230986565351486206e-01,2.360582351684570312e-01,1.008645594120025635e-01,7.829221338033676147e-02,3.777771070599555969e-02,-7.216563820838928223e-02,-1.401275862008333206e-03,-2.047472745180130005e-01,6.777143478393554688e-02,-6.283181905746459961e-02,6.008901819586753845e-02,1.078681647777557373e-02,-8.292602747678756714e-02,9.508222341537475586e-02,-3.038052320480346680e-01,-9.282774291932582855e-03,-3.551865741610527039e-02,1.192635446786880493e-01,2.436694316565990448e-02,-1.029372140765190125e-01,-6.831634789705276489e-02,-1.561976075172424316e-01,1.616667062044143677e-01,1.196196302771568298e-01,3.550394997000694275e-02,1.044736951589584351e-01,-2.743688225746154785e-02,-2.899760007858276367e-02,-1.935134828090667725e-02,-5.975026264786720276e-02,-2.912709861993789673e-02,7.869771867990493774e-02,-2.081265300512313843e-02,2.545703649520874023e-01,-3.451972082257270813e-02,2.073529548943042755e-02,1.078583225607872009e-01,-7.878972589969635010e-02,6.735565513372421265e-02,-1.186495944857597351e-01,-1.857072561979293823e-01,3.165216371417045593e-02,-1.029088348150253296e-01,9.516184777021408081e-02,1.370947808027267456e-02,7.616059482097625732e-02,5.157251656055450439e-02,2.565068937838077545e-02,3.097316250205039978e-02,-9.085205197334289551e-02,5.499069020152091980e-02,1.155302897095680237e-01,-1.005818322300910950e-02,-1.295643597841262817e-01,5.165000632405281067e-02,-6.884622573852539062e-02,-4.781063273549079895e-02,1.471960544586181641e-01,4.383899644017219543e-02,2.969204783439636230e-01,-2.518545649945735931e-02,-9.503652155399322510e-02,-1.449114363640546799e-02,1.703610718250274658e-01,-1.971014142036437988e-01,8.519279956817626953e-02,7.349193841218948364e-02,-2.027592808008193970e-01,9.589438326656818390e-03,-1.355729997158050537e-01,-1.144947297871112823e-02,3.680001199245452881e-02,-2.324504405260086060e-02,-1.736451667966321111e-04,-1.075484752655029297e-01,1.892208456993103027e-01,2.056821808218955994e-02,7.803399115800857544e-02,5.113979429006576538e-02,2.334306240081787109e-01,2.929230928421020508e-01,3.472810387611389160e-01,-9.320312179625034332e-03,-7.366197556257247925e-02,1.692025214433670044e-01,-1.445765141397714615e-02,5.596570968627929688e-01,2.679021656513214111e-01,5.611830390989780426e-03,-2.960789799690246582e-01,2.991384565830230713e-01,-1.749741286039352417e-01,-6.645976305007934570e-01,6.740671396255493164e-01,5.110760331153869629e-01,-1.659665405750274658e-01,-2.642334066331386566e-02,-2.859971225261688232e-01,-4.568833112716674805e-02,1.431521177291870117e-01,-5.061027780175209045e-02,2.677977383136749268e-01,3.864986076951026917e-02,8.352752029895782471e-02,2.676878571510314941e-01,-1.447378098964691162e-02,2.395460307598114014e-01,-3.265434131026268005e-02,-1.814712882041931152e-01,-4.817123711109161377e-02,-7.397264242172241211e-02,1.518321484327316284e-01,1.074417009949684143e-01,-6.164182722568511963e-02,1.080936193466186523e-01,-8.826810866594314575e-03,-1.271417886018753052e-01,9.689545631408691406e-02,-5.715501680970191956e-02,1.438101381063461304e-01,9.942378103733062744e-02,3.458409383893013000e-02,-5.431279912590980530e-02,-8.305248618125915527e-02,1.307578831911087036e-01,6.722307950258255005e-02,-8.878596872091293335e-02,1.486973911523818970e-01,-1.862957775592803955e-01,-1.011491864919662476e-01,-8.082222938537597656e-02,7.945100218057632446e-02,-1.447963565587997437e-01,1.374536305665969849e-01,1.353113949298858643e-01,-1.997535526752471924e-01,-1.447992622852325439e-01,2.581047639250755310e-02,-1.256135851144790649e-01,5.720512196421623230e-02,-1.750693470239639282e-01,1.461026258766651154e-02,9.184745699167251587e-02,-9.425931423902511597e-02,5.175523459911346436e-02,9.235849231481552124e-02,1.926688998937606812e-01,6.078736111521720886e-02,9.316221624612808228e-02,-6.492676585912704468e-02,2.445093728601932526e-02,6.090589985251426697e-02,1.612708717584609985e-02,-6.934259831905364990e-02,5.059774219989776611e-02,-3.425702452659606934e-02,1.663166582584381104e-01,-1.130852922797203064e-01,1.670292466878890991e-01,2.047598361968994141e-01,-4.387252405285835266e-02,-1.727919429540634155e-01,3.648624196648597717e-02,1.147893965244293213e-01,-1.129271686077117920e-01,-7.989731431007385254e-02,3.686897456645965576e-02,-6.191245838999748230e-02,1.059590578079223633e-01,3.332957625389099121e-01,1.263491660356521606e-01,8.616466075181961060e-02,1.578808426856994629e-01,-2.573181986808776855e-01,2.054274529218673706e-01,-1.985169351100921631e-01,-1.716416031122207642e-01,-6.487599015235900879e-02,1.683197319507598877e-01,-6.784933805465698242e-02,1.498868316411972046e-01,1.214449554681777954e-01,-2.278462052345275879e-02,-1.722159236669540405e-02,1.655252724885940552e-01,-5.820450186729431152e-02,-2.021321803331375122e-01,1.389960795640945435e-01,-2.438439615070819855e-02,3.680733963847160339e-02,1.567952521145343781e-02,-3.654563054442405701e-02,-8.595662564039230347e-02,7.368671149015426636e-02,2.080126553773880005e-01,-5.656849220395088196e-02,-5.537661910057067871e-02,-5.598208308219909668e-02,2.033397108316421509e-01,6.031342968344688416e-02,-1.445585489273071289e-02,-8.706968277692794800e-03,1.569439657032489777e-02,1.321733146905899048e-01,5.780521035194396973e-02,-1.110171452164649963e-01,3.894703686237335205e-01,-1.812738478183746338e-01,2.283367216587066650e-01,7.021525874733924866e-03,3.376605212688446045e-01,1.192678883671760559e-02,-7.637096643447875977e-01,1.151919830590486526e-02,3.825847506523132324e-01,-1.199142038822174072e-01,1.597879640758037567e-02,-4.512070119380950928e-02,-4.136779606342315674e-01,-2.322103083133697510e-01,9.655947238206863403e-02,1.030356856063008308e-03,-2.644611001014709473e-01,-2.742321193218231201e-01,1.568390876054763794e-01,1.087251752614974976e-01,1.253557801246643066e-01,2.499288134276866913e-02,1.186901256442070007e-01,4.775649681687355042e-02,1.578856259584426880e-01,1.751341521739959717e-01,2.628433108329772949e-01,2.662527263164520264e-01,2.071907073259353638e-01,-1.029616072773933411e-01,2.003372311592102051e-01,1.374835819005966187e-01,1.230700984597206116e-01,1.524515599012374878e-01,2.420096248388290405e-01,1.459203753620386124e-02,1.397923082113265991e-01,-2.562743052840232849e-02,1.644181758165359497e-01,2.223161607980728149e-01,4.724684357643127441e-02,-2.508093416690826416e-01,-3.685732558369636536e-02,-8.177562057971954346e-02,1.173208951950073242e-01,-1.467597633600234985e-01,2.405925840139389038e-01,2.120443247258663177e-02,-2.268977612257003784e-01,2.832765579223632812e-01,-2.502555549144744873e-01,1.340543329715728760e-01,-7.268548943102359772e-03,-2.514312267303466797e-01,-9.737252444028854370e-02,-1.851898990571498871e-02,-2.758130133152008057e-01,-1.493088901042938232e-01,-1.940908841788768768e-02,-1.084841862320899963e-01,1.717299669981002808e-01,-1.494039595127105713e-01,2.383804619312286377e-01,-1.988504379987716675e-01,6.095692515373229980e-02,-3.051739372313022614e-02,3.736748099327087402e-01,1.452666819095611572e-01,9.182056039571762085e-02,2.844219803810119629e-01,-3.169150948524475098e-01,5.016106367111206055e-01,2.166341394186019897e-01,2.477407082915306091e-02,9.800371527671813965e-02,2.073259800672531128e-01,-3.669050056487321854e-03,-3.649210184812545776e-02,-9.195020049810409546e-02,-1.088774353265762329e-01,1.236683428287506104e-01,1.197806559503078461e-02,-3.207577392458915710e-02,-2.513998001813888550e-02,-1.392220258712768555e-01,-7.117275893688201904e-02,-4.719172418117523193e-02,-3.651745319366455078e-01,1.016260012984275818e-01,-2.066573053598403931e-01,-1.179236248135566711e-01,4.454509541392326355e-02,-1.994255334138870239e-01,-2.474335208535194397e-02,-1.157272979617118835e-01,1.311783641576766968e-01,-1.484084315598011017e-02,2.213118970394134521e-01,1.751638203859329224e-02,-9.321501106023788452e-02,1.531160771846771240e-01,1.906989887356758118e-02,7.707899808883666992e-02,2.758827209472656250e-01,-7.586433552205562592e-03,-5.082147940993309021e-02,-3.325645998120307922e-02,-3.494461998343467712e-02,2.462530136108398438e-02,1.179282069206237793e-01,3.266915977001190186e-01,-2.081049978733062744e-02,-6.272995471954345703e-02,1.661009192466735840e-01,1.732306331396102905e-01,2.158563137054443359e-01,6.514336168766021729e-02,4.085751995444297791e-02,1.216489821672439575e-01,1.701028943061828613e-01,-2.824357748031616211e-01,1.562914401292800903e-01,2.640362977981567383e-01,8.865283429622650146e-02,8.734606951475143433e-02,1.268353164196014404e-01,1.491427570581436157e-01,8.871096372604370117e-02,5.303507670760154724e-02,1.551600396633148193e-01,1.710316240787506104e-01,1.624363064765930176e-01,-1.988599002361297607e-01,-2.644401192665100098e-01,1.402551680803298950e-01,5.557774752378463745e-02,-3.510542213916778564e-01,-3.792574405670166016e-01,4.700138047337532043e-02,5.085975397378206253e-03,3.252378478646278381e-02,4.250177741050720215e-01,3.423853591084480286e-02,-4.960802793502807617e-01,1.628195643424987793e-01,-8.236531168222427368e-02,-6.157244443893432617e-01,2.398778498172760010e-01,1.766877919435501099e-01,-2.274876646697521210e-02,-5.242252256721258163e-03,-1.694621518254280090e-02,5.678001418709754944e-02,1.138336360454559326e-01,-8.943605422973632812e-02,8.793036639690399170e-02,1.320666372776031494e-01,-3.954850509762763977e-02,-2.547992393374443054e-02,3.555523604154586792e-02,1.907197684049606323e-01,-1.012812554836273193e-01,-4.020179435610771179e-02,1.481265295296907425e-02,-9.051078557968139648e-02,1.360332667827606201e-01,9.136970341205596924e-02,8.061093837022781372e-02,-3.110872814431786537e-03,-1.966172270476818085e-02,-1.442643260816112161e-04,4.223778843879699707e-02,3.656769171357154846e-02,1.189208496361970901e-02,1.237192824482917786e-01,-2.078293822705745697e-03,-8.341279812157154083e-03,1.161844730377197266e-01,7.006292045116424561e-02,2.654969394207000732e-01,3.099929988384246826e-01,-6.713202595710754395e-02,-4.953456670045852661e-02,8.231014758348464966e-02,-2.862262427806854248e-01,1.256072148680686951e-02,-7.204607874155044556e-02,8.200196549296379089e-03,-1.929907687008380890e-02,1.796789467334747314e-02,6.726364046335220337e-02,-8.521347492933273315e-02,-1.339051127433776855e-01,6.471113860607147217e-02,2.133182995021343231e-02,1.184187084436416626e-01,-1.094449982047080994e-01,-1.902303695678710938e-01,-4.929348453879356384e-02,3.059969842433929443e-02,7.797027379274368286e-02,1.326819509267807007e-01,-1.452069729566574097e-01,-2.013838738203048706e-01,9.135934710502624512e-02,8.741638809442520142e-02,-5.721065029501914978e-02,-6.497509777545928955e-02,-7.909812033176422119e-02,-2.262309193611145020e-02,-1.132673025131225586e-01,1.981829851865768433e-01,-1.001199856400489807e-01,-2.943236846476793289e-03,4.170941188931465149e-02,-1.185101270675659180e-01,1.282952725887298584e-01,-9.613715857267379761e-02,-1.489401161670684814e-01,4.341379553079605103e-02,-1.282791942358016968e-01,-1.449230909347534180e-01,-3.206847235560417175e-02,-2.047597058117389679e-02,-3.803251544013619423e-03,-2.211529389023780823e-02,8.222504705190658569e-02,-1.909977197647094727e-01,-6.378269940614700317e-02,-1.305363029241561890e-01,-1.957147866487503052e-01,2.440135926008224487e-02,-1.481731142848730087e-02,1.940115913748741150e-02,7.732482254505157471e-02,-3.290917724370956421e-02,1.341988332569599152e-02,9.457019716501235962e-02,1.177925802767276764e-02,2.265624236315488815e-03,-2.234340086579322815e-02,8.195963688194751740e-03,-4.220542311668395996e-02,8.144910633563995361e-02,-1.506609022617340088e-01,1.611797660589218140e-01,1.833299845457077026e-01,-1.314008086919784546e-01,-7.299738377332687378e-02,6.732426583766937256e-02,1.849891692399978638e-01,-7.176375389099121094e-02,5.660580936819314957e-03,-4.195747897028923035e-02,-3.490515798330307007e-02,5.809704586863517761e-02,1.239352021366357803e-02,2.441540360450744629e-02,4.727337062358856201e-01,-9.526423215866088867e-01,-9.683986902236938477e-01,1.115965366363525391e+00,5.622525215148925781e-01,-8.489467501640319824e-01,2.523935437202453613e-01,2.379070967435836792e-01,6.706213206052780151e-02,3.464241325855255127e-01,1.292799860239028931e-01,-2.150530554354190826e-02,-8.036924600601196289e-01,-9.874364137649536133e-01,-4.972656071186065674e-01,-1.576442122459411621e-01,1.527972221374511719e-01,2.082870900630950928e-01,2.494367212057113647e-01,-1.240093410015106201e-01,1.148297451436519623e-02,-1.099322289228439331e-01,-9.023674577474594116e-02,1.695354580879211426e-01,1.599134877324104309e-03,1.359329372644424438e-01,5.774929001927375793e-02,8.727262169122695923e-02,2.995097637176513672e-02,1.397419422864913940e-01,2.511543780565261841e-02,6.238651648163795471e-02,2.156476825475692749e-01,2.116920202970504761e-01,1.783205419778823853e-01,1.288940012454986572e-01,2.549798488616943359e-01,-1.208158093504607677e-03,-1.214666888117790222e-01,3.740962445735931396e-01,-3.119483962655067444e-02,1.397333443164825439e-01,1.074238792061805725e-01,8.345821499824523926e-02,3.776837885379791260e-01,7.747357338666915894e-02,-5.038021132349967957e-02,5.148956775665283203e-01,1.408054232597351074e-01,-1.150845661759376526e-01,1.330581214278936386e-02,5.118693411350250244e-02,4.559218510985374451e-02,-1.835397183895111084e-01,7.072634994983673096e-02,9.008940309286117554e-02,1.141012459993362427e-01,-2.389682382345199585e-01,1.368290930986404419e-01,-1.775007247924804688e-01,-2.060741484165191650e-01,-1.267988830804824829e-01,1.727024912834167480e-01,2.108477950096130371e-01,-1.646388471126556396e-01,-2.511967420578002930e-01,7.017033174633979797e-03,2.791520655155181885e-01,6.212844979017972946e-03,8.079923689365386963e-02,6.541586667299270630e-02,2.007054984569549561e-01,2.596695423126220703e-01,-4.336170107126235962e-02,2.770919501781463623e-01,-1.013183221220970154e-01,-8.592540025711059570e-02,-1.894620507955551147e-01,-2.286358028650283813e-01,1.609836369752883911e-01,-2.648130357265472412e-01,-4.578446447849273682e-01,5.552702397108078003e-02,2.865148521959781647e-02,-1.732976287603378296e-01,1.168414130806922913e-01,-2.266460061073303223e-01,4.435078799724578857e-02,-1.236633118242025375e-02,-2.374881356954574585e-01,2.077378183603286743e-01,-1.003839001059532166e-01,-2.959598600864410400e-01,7.650348823517560959e-03,1.046140342950820923e-01,3.201979994773864746e-01,-6.568681565113365650e-04,3.545404970645904541e-01,2.926314175128936768e-01,-9.080765396356582642e-02,6.576602905988693237e-02,2.160100191831588745e-01,9.833301603794097900e-02,-1.411784905940294266e-02,-1.065702214837074280e-01,2.169614424929022789e-03,2.872113883495330811e-02,1.885773688554763794e-01,-5.420678481459617615e-02,6.588017940521240234e-02,2.129836706444621086e-03,2.732092738151550293e-01,1.278383731842041016e-01,-1.286749690771102905e-01,4.921238124370574951e-02,1.572323888540267944e-01,-1.047752797603607178e-01,1.055460125207901001e-01,-1.283281743526458740e-01,-4.203576967120170593e-02,3.465801849961280823e-02,6.188576668500900269e-02,-1.179015822708606720e-02,-1.860799938440322876e-01,8.331302087754011154e-04,2.024499624967575073e-01,3.626270592212677002e-01,5.192021727561950684e-01,5.100845098495483398e-01,2.272012084722518921e-01,-2.226626425981521606e-01,-4.689000844955444336e-01,-1.839854866266250610e-01,9.739734232425689697e-02,4.703223705291748047e-01,9.088392555713653564e-02,1.500865910202264786e-02,9.809152036905288696e-02,1.510337889194488525e-01,-1.934976899065077305e-03,-2.264406383037567139e-01,-6.487185955047607422e-01,-8.378006815910339355e-01,-7.971260547637939453e-01,-4.954192638397216797e-01,-2.713887989521026611e-01,-3.512001037597656250e-01,-6.244751214981079102e-01,-4.393753707408905029e-01,-5.759497284889221191e-01,-2.332922667264938354e-01,-3.836019337177276611e-01,-2.353938370943069458e-01,-3.125010728836059570e-01,-8.533917367458343506e-02,-2.152969837188720703e-01,7.955909520387649536e-02,8.951836824417114258e-02,-1.007588133215904236e-01,-8.201099932193756104e-02,1.277243345975875854e-01,-4.569659940898418427e-03,-2.331376634538173676e-02,1.747729023918509483e-03,2.013573646545410156e-01,1.881647706031799316e-01,6.111001595854759216e-02,1.763990670442581177e-01,2.019171118736267090e-01,3.010985553264617920e-01,1.852870285511016846e-01,2.064862102270126343e-01,2.511513531208038330e-01,2.347905039787292480e-01,2.153710871934890747e-01,-4.725488834083080292e-03,9.288479387760162354e-02,-1.145128458738327026e-01,8.985693007707595825e-02,1.892805993556976318e-01,9.802240878343582153e-02,1.159583032131195068e-01,4.810172691941261292e-02,2.263849601149559021e-02,-7.031312584877014160e-02,-9.780356287956237793e-02,8.087783306837081909e-02,-1.809016317129135132e-01,-3.874167799949645996e-02,7.943062111735343933e-03,-6.573629379272460938e-02,6.803462654352188110e-02,-9.915065020322799683e-02,1.012928485870361328e-01,-1.226266026496887207e-01,1.412642896175384521e-01,9.038345515727996826e-02,1.883030310273170471e-02,1.314334422349929810e-01,-2.188625745475292206e-02,2.940866537392139435e-02,6.256588734686374664e-03,8.934940211474895477e-03,1.915486305952072144e-01,1.973392367362976074e-01,1.486583650112152100e-01,2.609265595674514771e-02,-3.776717232540249825e-03,-9.418852627277374268e-03,1.613480746746063232e-01,2.770119011402130127e-01,7.042096555233001709e-02,1.279187798500061035e-01,2.037594467401504517e-01,-9.808833710849285126e-03,1.179930344223976135e-01,-4.373666644096374512e-02,2.651540637016296387e-01,1.004228591918945312e-01,1.608752310276031494e-01,1.321744769811630249e-01,1.785648018121719360e-01,2.263544350862503052e-01,1.426501572132110596e-01,-2.082459442317485809e-02,4.371062815189361572e-01,1.530244108289480209e-02,2.870449721813201904e-01,1.804132908582687378e-01,5.178901553153991699e-02,3.522001802921295166e-01,6.051355227828025818e-02,1.769441813230514526e-01,8.951232582330703735e-02,2.882507443428039551e-02,4.481187462806701660e-02,2.240322530269622803e-01,1.066040843725204468e-01,1.620966196060180664e-02,1.868079900741577148e-01,-8.357720077037811279e-02,-6.907959282398223877e-02,2.583028189837932587e-02,-1.109675690531730652e-02,8.006370626389980316e-03,7.238563895225524902e-02,2.297206036746501923e-02,1.228331178426742554e-01,2.436908707022666931e-02,1.237533017992973328e-01,1.117848232388496399e-01,1.666666567325592041e-01,-1.057550497353076935e-02,2.218678742647171021e-01,2.079626321792602539e-01,5.827291011810302734e-01,6.852402687072753906e-01,4.226052463054656982e-01,3.039394319057464600e-01,2.459927201271057129e-01,3.956699073314666748e-01,4.288652837276458740e-01,-1.199669986963272095e-01,4.553144872188568115e-01,1.962838321924209595e-01,-2.421817928552627563e-01,6.956008076667785645e-02,-1.890045404434204102e-01,1.639902358874678612e-03,4.036978781223297119e-01,1.484436988830566406e-01,1.665644496679306030e-01,1.137938126921653748e-01,-1.966261863708496094e-01,5.148333311080932617e-02,-2.417005747556686401e-01,-1.602289080619812012e-01,8.443330228328704834e-02,-1.976093947887420654e-01,1.438007876276969910e-02,-6.142470613121986389e-02,-1.420667320489883423e-01,-5.861635878682136536e-02,-1.593414247035980225e-01,1.880273409187793732e-02,-9.998465888202190399e-03,3.554236516356468201e-02,7.925789058208465576e-02,-1.319591188803315163e-03,-1.246945858001708984e-01,1.134144067764282227e-01,-5.778913944959640503e-02,1.204620972275733948e-01,1.036474332213401794e-01,2.241288572549819946e-01,-2.884369902312755585e-02,2.872578799724578857e-01,-4.555732756853103638e-02,2.225508987903594971e-01,-7.160489261150360107e-02,-2.948704920709133148e-02,4.265005514025688171e-02,5.147395282983779907e-02,-1.248668581247329712e-01,3.780346363782882690e-02,-7.529974728822708130e-02,1.726603694260120392e-02,1.304767727851867676e-01,1.949221938848495483e-01,-1.138305291533470154e-02,1.283098012208938599e-01,1.049685180187225342e-01,-1.377262920141220093e-01,2.058669477701187134e-01,1.132107712328433990e-02,4.257582500576972961e-02,-1.430011093616485596e-01,9.689304046332836151e-03,-1.525093466043472290e-01,-5.850138142704963684e-02,-1.769078969955444336e-01,5.638798698782920837e-03,1.222907006740570068e-01,-5.411321297287940979e-02,-7.249010354280471802e-02,-9.903898835182189941e-02,-5.687761679291725159e-02,-2.747875154018402100e-01,-6.800738722085952759e-02,-3.450696766376495361e-01,-9.073706343770027161e-03,8.299160748720169067e-02,1.678718328475952148e-01,9.125961363315582275e-02,-1.653965860605239868e-01,2.880944609642028809e-01,-1.751377284526824951e-01,-8.920015394687652588e-02,2.057643383741378784e-01,5.638929083943367004e-02,9.047846309840679169e-03,-2.394968271255493164e-02,-1.394613683223724365e-01,4.401495307683944702e-02,5.335658416152000427e-02,-4.726697877049446106e-02,5.525279417634010315e-02,-6.052866578102111816e-02,1.633741110563278198e-01,2.245084941387176514e-02,7.462608814239501953e-02,-8.563823997974395752e-02,-8.827047795057296753e-02,2.007955312728881836e-01,-5.125345289707183838e-02,1.083375234156847000e-02,-9.963083267211914062e-02,-1.234357431530952454e-01,-7.055723667144775391e-02,1.904234886169433594e-01,5.887345224618911743e-02,5.362937226891517639e-02,-1.281675547361373901e-01,5.911789089441299438e-02,-2.703308127820491791e-03,-4.645418841391801834e-03,-5.582652986049652100e-02,1.156948693096637726e-02,-1.124745011329650879e-01,-1.672277040779590607e-02,-5.338333174586296082e-02,4.395567812025547028e-03,-3.385889530181884766e-02,-4.035931080579757690e-02,1.200505346059799194e-01,-1.486072391271591187e-01,1.427377760410308838e-01,4.661733657121658325e-02,2.830590605735778809e-01,1.668400913476943970e-01,8.314250409603118896e-02,1.387589424848556519e-01,7.896072417497634888e-02,1.255486309528350830e-01,3.823397755622863770e-01,1.919494569301605225e-01,4.133200049400329590e-01,9.015380591154098511e-02,-2.556116878986358643e-01,1.092869937419891357e-01,-1.947639286518096924e-01,4.527266025543212891e-01,6.070288270711898804e-02,-2.584054693579673767e-02,1.298940181732177734e-01,2.822883129119873047e-01,7.613944411277770996e-01,6.288247108459472656e-01,6.679862737655639648e-01,4.286323189735412598e-01,7.258780598640441895e-01,7.191877961158752441e-01,9.788619279861450195e-01,6.356813907623291016e-01,6.647245883941650391e-01,7.522597312927246094e-01,4.086832404136657715e-01,5.869017243385314941e-01,4.059696495532989502e-01,1.313670575618743896e-01,4.669856131076812744e-01,2.370035350322723389e-01,2.243708819150924683e-01,3.454623371362686157e-02,1.852635443210601807e-01,1.045350730419158936e-01,1.328025013208389282e-01,-1.134296879172325134e-01,-1.322030723094940186e-01,1.511588245630264282e-01,-2.789474278688430786e-02,5.805407185107469559e-03,-9.043869376182556152e-02,6.660116463899612427e-02,-2.173287570476531982e-01,-3.062795102596282959e-01,2.649064362049102783e-02,-1.793597042560577393e-01,1.538276970386505127e-01,-2.193829864263534546e-01,1.923917531967163086e-01,-1.765129566192626953e-01,1.734465956687927246e-01,1.911193281412124634e-01,2.755689993500709534e-02,9.396158903837203979e-02,4.623237252235412598e-02,-1.250826567411422729e-01,9.910140186548233032e-02,-1.699882373213768005e-02,-1.655747741460800171e-01,9.622088074684143066e-02,-8.520791679620742798e-02,-2.879169397056102753e-02,1.487938910722732544e-01,-1.641035526990890503e-01,-5.060535669326782227e-02,2.374791502952575684e-01,2.640470862388610840e-01,4.517933353781700134e-03,1.980386525392532349e-01,1.077273041009902954e-01,-2.966157719492912292e-02,-1.579282805323600769e-02,1.006059721112251282e-01,3.207172267138957977e-03,2.596196532249450684e-01,4.713086038827896118e-02,3.371104598045349121e-01,9.841845929622650146e-02,1.823777705430984497e-01,-2.198508530855178833e-01,1.709640622138977051e-01,-3.576312959194183350e-01,4.904023557901382446e-02,-1.888312697410583496e-01,3.938145190477371216e-02,1.594133824110031128e-01,-4.966327548027038574e-02,-1.017902884632349014e-02,1.113322451710700989e-01,-8.712708204984664917e-02,-1.258390992879867554e-01,-5.174351111054420471e-02,-4.127714782953262329e-02,-8.574488013982772827e-02,-1.326052397489547729e-01,2.906209044158458710e-02,-2.585966885089874268e-01,-4.851242527365684509e-03,-2.959745526313781738e-01,-3.111799061298370361e-01,-1.185666471719741821e-01,-1.783578470349311829e-02,-1.330411732196807861e-01,-1.444811373949050903e-01,-3.026174306869506836e-01,1.130181029438972473e-01,-2.768821120262145996e-01,-8.701410889625549316e-02,-2.049572318792343140e-01,-3.081521093845367432e-01,-4.798658192157745361e-03,1.529962569475173950e-01,-1.990439146757125854e-01,-2.170781940221786499e-01,2.206964492797851562e-01,-8.977482467889785767e-02,-2.195162624120712280e-01,-1.137224957346916199e-01,-1.114687845110893250e-01,-4.124783724546432495e-02,-2.054465711116790771e-01,4.653508961200714111e-02,-1.580305397510528564e-01,9.223969280719757080e-02,-5.026848316192626953e-01,-1.020480021834373474e-01,1.180650144815444946e-01,-4.211431443691253662e-01,-2.279297262430191040e-02,-1.792571395635604858e-01,-1.490917056798934937e-01,4.245139062404632568e-01,2.339401096105575562e-01,-1.371203809976577759e-01,1.335296686738729477e-02,-2.206559106707572937e-02,3.860106766223907471e-01,-7.895590662956237793e-01,3.101220428943634033e-01,3.410652875900268555e-01,2.310179620981216431e-01,1.944981515407562256e-01,1.007202193140983582e-01,4.593634605407714844e-02,1.558400988578796387e-01,2.004333883523941040e-01,9.816525131464004517e-02,3.349725604057312012e-01,2.563640773296356201e-01,2.191550880670547485e-01,1.889916807413101196e-01,1.669982224702835083e-01,1.157895475625991821e-01,1.975189745426177979e-01,1.748383194208145142e-01,3.593252301216125488e-01,2.586624324321746826e-01,1.559654176235198975e-01,2.995968796312808990e-02,1.358238607645034790e-01,1.597530841827392578e-01,6.129888072609901428e-02,1.287584751844406128e-01,-3.299800306558609009e-02,-1.041386425495147705e-01,2.087793350219726562e-01,2.964749000966548920e-02,2.906259596347808838e-01,1.693434715270996094e-01,5.086383968591690063e-02,9.093750268220901489e-02,-2.900868467986583710e-02,5.143247544765472412e-02,3.411704301834106445e-02,2.880310080945491791e-02,-7.947243750095367432e-02,1.833390295505523682e-01,-2.134713530540466309e-01,9.318259358406066895e-02,-1.882264390587806702e-02,-8.970747143030166626e-02,7.551503181457519531e-02,1.207311898469924927e-01,4.024701565504074097e-02,1.701105833053588867e-01,-1.919572204351425171e-01,3.802163153886795044e-02,1.659157425165176392e-01,2.249189466238021851e-01,1.699155867099761963e-01,7.529576122760772705e-02,4.465122148394584656e-02,-3.313054144382476807e-02,7.069668173789978027e-02,6.671275198459625244e-02,3.778479695320129395e-01,-3.359755128622055054e-02,2.882138788700103760e-01,7.812269777059555054e-02,-1.422116011381149292e-01,1.633932888507843018e-01,7.191594690084457397e-02,-3.087279200553894043e-01,-9.609597921371459961e-02,9.948955848813056946e-03,9.889889508485794067e-02,2.531620264053344727e-01,-1.484955549240112305e-01,4.883767291903495789e-02,-5.278110504150390625e-02,-2.697815895080566406e-01,1.357145309448242188e-01,-1.727140694856643677e-01,1.464380770921707153e-01,-1.486711110919713974e-02,-5.727973207831382751e-02,-2.786490619182586670e-01,2.543626129627227783e-01,6.190706416964530945e-02,-3.193286955356597900e-01,-2.991230785846710205e-02,-4.169974625110626221e-01,6.639435887336730957e-02,7.148016244173049927e-02,-4.335653036832809448e-03,-8.797799795866012573e-02,1.682624816894531250e-01,1.813124120235443115e-01,-1.430575251579284668e-01,1.721735447645187378e-01,-9.921076893806457520e-02,-1.645226627588272095e-01,7.081935554742813110e-02,5.636121705174446106e-02,7.704451680183410645e-03,-4.480496421456336975e-02,-2.973631583154201508e-02,-1.261681504547595978e-02,1.442302018404006958e-01,1.864746958017349243e-01,1.291276216506958008e-01,1.217148602008819580e-01,-1.689191907644271851e-01,5.928743630647659302e-02,4.401450231671333313e-02,1.308848708868026733e-01,1.154345422983169556e-01,-1.804474145174026489e-01,-6.958601623773574829e-02,2.548460364341735840e-01,2.042754739522933960e-01,1.615671813488006592e-01,1.406262964010238647e-01,-2.845165431499481201e-01,-1.518948972225189209e-01,-1.611388325691223145e-01,-2.737249135971069336e-01,-2.621858417987823486e-01,-1.730663925409317017e-01,-4.377865195274353027e-01,-5.062648057937622070e-01,2.349456772208213806e-02,1.434291750192642212e-01,8.330332040786743164e-01,7.694554328918457031e-01,4.948168694972991943e-01,-7.180818915367126465e-02,1.472966372966766357e-01,3.958906829357147217e-01,-2.830893397331237793e-01,-6.801868677139282227e-01,1.559848785400390625e-01,1.753408163785934448e-01,1.888591647148132324e-01,4.999693930149078369e-01,2.713595628738403320e-01,1.687965840101242065e-01,-7.050364464521408081e-02,-7.635032385587692261e-02,-2.535781860351562500e-01,-4.773127846419811249e-03,1.519059091806411743e-01,-3.639306128025054932e-02,7.613504678010940552e-02,-7.876231521368026733e-02,1.106265261769294739e-01,3.653056919574737549e-01,-7.969317585229873657e-02,4.023301973938941956e-02,-2.952444832772016525e-03,-1.887849718332290649e-02,-6.444857455790042877e-03,6.224972382187843323e-02,8.746765553951263428e-02,-1.313134282827377319e-01,8.924893289804458618e-02,1.307076541706919670e-03,1.489989906549453735e-01,-4.116903245449066162e-02,1.901100575923919678e-01,2.290278971195220947e-01,-1.551095694303512573e-01,1.412630379199981689e-01,3.987379744648933411e-02,-1.739287227392196655e-01,-1.273187845945358276e-01,-9.384039789438247681e-02,-2.132421135902404785e-01,-1.031102053821086884e-02,1.893593817949295044e-01,-2.613190747797489166e-02,7.197244465351104736e-02,1.454360187053680420e-01,-1.777701079845428467e-01,-2.270150631666183472e-01,-1.237686350941658020e-01,1.840328797698020935e-02,-1.775733381509780884e-01,2.367413341999053955e-01,-1.910639107227325439e-01,4.417350888252258301e-02,-2.282558530569076538e-01,-1.476555317640304565e-01,-2.014051079750061035e-01,-4.917169362306594849e-02,-1.317082643508911133e-01,-1.226217523217201233e-01,1.069581955671310425e-01,-1.021934300661087036e-01,1.415889263153076172e-01,-2.118941992521286011e-01,6.283421814441680908e-02,2.902026772499084473e-01,2.642525732517242432e-01,-1.327590197324752808e-01,1.784160584211349487e-01,-3.885817527770996094e-02,1.132667139172554016e-01,4.932921845465898514e-03,-6.187309697270393372e-02,3.173714280128479004e-01,-4.101642668247222900e-01,-2.113666385412216187e-02,-7.824723422527313232e-02,7.988887280225753784e-02,-4.141466319561004639e-02,-9.470642544329166412e-03,-7.976195961236953735e-02,1.369839906692504883e-01,-4.751781225204467773e-01,-6.981372833251953125e-02,-4.631811007857322693e-02,-6.931539624929428101e-02,-3.340736776590347290e-02,1.026161685585975647e-01,2.224273420870304108e-02,2.072398662567138672e-01,3.616756875999271870e-04,-2.587908208370208740e-01,7.599691301584243774e-02,-8.184539526700973511e-02,3.398785740137100220e-02,-2.672413289546966553e-01,-9.692870825529098511e-02,6.925562769174575806e-02,6.027085706591606140e-03,-1.619971394538879395e-01,2.116417288780212402e-01,2.609548531472682953e-02,1.671373397111892700e-01,-5.509947240352630615e-02,-7.711293548345565796e-02,9.211045503616333008e-02,1.331427544355392456e-01,-1.372023373842239380e-01,-1.799138337373733521e-01,2.476003393530845642e-02,2.062282711267471313e-02,1.545435488224029541e-01,3.192920088768005371e-01,-2.994341552257537842e-01,2.931767404079437256e-01,6.782887876033782959e-02,1.314813643693923950e-01,-1.149998977780342102e-01,-1.841798573732376099e-01,-4.411765336990356445e-01,-6.757512092590332031e-01,4.207124933600425720e-03,5.304787158966064453e-01,2.129307389259338379e-01,-1.006492227315902710e-01,-2.378382682800292969e-01,4.919681549072265625e-01,5.405007302761077881e-02,9.750638157129287720e-03,1.388392597436904907e-01,-1.884981058537960052e-02,-1.928160488605499268e-01,7.299953103065490723e-01,2.199220508337020874e-01,-2.050085216760635376e-01,5.006049945950508118e-02,-1.421987451612949371e-02,-3.744550421833992004e-02,-3.898786148056387901e-03,5.495267733931541443e-02,-1.440359055995941162e-01,1.755570806562900543e-02,2.042363863438367844e-03,-1.536547094583511353e-01,4.874577373266220093e-02,-7.426231354475021362e-02,2.446755394339561462e-02,-3.820474073290824890e-02,-1.280339807271957397e-01,-4.546315595507621765e-02,-2.842151373624801636e-02,8.246731013059616089e-02,-2.472190931439399719e-02,-4.508957266807556152e-02,-3.487443923950195312e-02,1.117029264569282532e-01,4.372176155447959900e-02,7.840679585933685303e-02,-2.409858070313930511e-02,6.163920834660530090e-02,1.149429604411125183e-01,7.065568864345550537e-02,2.385822823271155357e-03,1.228253617882728577e-01,1.277848146855831146e-02,8.435490727424621582e-02,8.590666949748992920e-02,-5.112435296177864075e-02,-7.118750363588333130e-02,1.689439564943313599e-01,-3.474541008472442627e-02,-3.755690529942512512e-02,-3.929460793733596802e-02,-6.234410777688026428e-02,1.234380714595317841e-02,-3.242244198918342590e-02,4.238623194396495819e-03,-7.616367936134338379e-02,2.991056069731712341e-02,-8.028412610292434692e-02,1.789462417364120483e-01,-1.868812716566026211e-03,-4.146562423557043076e-03,-5.486308783292770386e-02,5.535012111067771912e-02,-1.258019506931304932e-01,-7.855030894279479980e-02,-3.416979312896728516e-02,-1.246717050671577454e-01,1.773130446672439575e-01,-1.664438545703887939e-01,4.921010136604309082e-02,-2.267074398696422577e-02,-9.397853910923004150e-02,5.072906496934592724e-04,9.394113905727863312e-03,-1.466102898120880127e-01,1.514739543199539185e-01,-1.655934453010559082e-01,1.612128913402557373e-01,-3.127655247226357460e-03,-4.558479413390159607e-02,1.206555441021919250e-01,4.191228374838829041e-02,-1.454896032810211182e-01,1.752282492816448212e-02,-1.165452376008033752e-01,-5.023838952183723450e-02,-7.274807244539260864e-02,-2.806889638304710388e-02,2.812261134386062622e-02,-2.344900518655776978e-01,4.761604592204093933e-02,-1.434403657913208008e-01,3.359604999423027039e-02,-2.155888080596923828e-01,-1.028171405196189880e-01,-9.240641444921493530e-02,-9.934887290000915527e-03,-1.025201473385095596e-02,-6.856817007064819336e-02,-3.876260295510292053e-02,-1.636468172073364258e-01,-5.715657025575637817e-02,-6.433968245983123779e-02,-1.341775357723236084e-01,7.666137814521789551e-02,-5.925538763403892517e-02,2.404562430456280708e-03,-2.109723538160324097e-01,2.590204775333404541e-02,-7.831685245037078857e-02,-1.103839650750160217e-01,7.154628634452819824e-02,-9.224347025156021118e-02,-8.757005445659160614e-03,3.320028632879257202e-02,-8.994955569505691528e-03,-1.138165146112442017e-01,9.013355523347854614e-02,-7.546217739582061768e-02,-1.742251217365264893e-01,2.927516996860504150e-01,-2.893903106451034546e-02,3.065226599574089050e-02,2.088810354471206665e-01,2.154102921485900879e-01,1.091030240058898926e-01,4.367803931236267090e-01,-4.452988505363464355e-01,-1.205657720565795898e+00,7.319428324699401855e-01,3.105916678905487061e-01,-8.503431081771850586e-02,1.822073906660079956e-01,4.421239793300628662e-01,-1.286063939332962036e-01,-2.013961970806121826e-01,3.086365461349487305e-01,4.893090426921844482e-01,5.086427330970764160e-01,3.968190550804138184e-01,2.576106190681457520e-01,2.514838576316833496e-01,2.930352091789245605e-01,1.339850127696990967e-01,3.856100887060165405e-02,-4.622703790664672852e-02,3.823471069335937500e-02,1.186072155833244324e-01,2.634907960891723633e-01,1.368056386709213257e-01,7.297031581401824951e-02,2.655484080314636230e-01,-1.557153016328811646e-01,2.918868362903594971e-01,2.045777291059494019e-01,6.644130498170852661e-02,3.871417045593261719e-01,1.367088705301284790e-01,1.714097708463668823e-01,1.192110106348991394e-01,8.301032334566116333e-02,1.643315702676773071e-01,1.607765108346939087e-01,2.172952145338058472e-01,8.616424351930618286e-02,5.219501256942749023e-02,-8.918390423059463501e-02,7.789735496044158936e-02,-5.007470957934856415e-03,4.342895001173019409e-02,8.180185407400131226e-02,7.064881734549999237e-03,-5.393844470381736755e-02,1.009424775838851929e-02,3.750009462237358093e-02,2.922598123550415039e-01,-2.013167589902877808e-01,2.324614375829696655e-01,1.434691995382308960e-01,1.030764654278755188e-01,2.404997497797012329e-01,2.242244221270084381e-02,1.195006221532821655e-01,2.396375536918640137e-01,2.111660838127136230e-01,2.229768335819244385e-01,7.441734522581100464e-02,1.573350466787815094e-02,1.493203490972518921e-01,1.106968894600868225e-01,4.937524199485778809e-01,2.675774395465850830e-01,-3.485628962516784668e-02,1.307782083749771118e-01,1.186861842870712280e-01,4.457398056983947754e-01,2.518717646598815918e-01,2.641805410385131836e-01,1.154934987425804138e-01,1.371820271015167236e-01,3.652333617210388184e-01,-2.832660377025604248e-01,-1.048004776239395142e-01,-9.833151847124099731e-02,7.636447995901107788e-02,1.675887256860733032e-01,-3.104854226112365723e-01,-4.781076312065124512e-02,-1.806190237402915955e-02,-3.255238831043243408e-01,-2.325187474489212036e-01,-1.065796911716461182e-01,-3.179083764553070068e-01,-4.920406267046928406e-02,-3.403505682945251465e-01,3.778834640979766846e-02,-1.245096549391746521e-01,-2.103211358189582825e-02,-2.000946253538131714e-01,-3.011123836040496826e-01,3.637712821364402771e-02,-2.883451581001281738e-01,5.784584581851959229e-02,-1.115496084094047546e-01,-3.487361129373311996e-03,1.138525605201721191e-01,-9.026136249303817749e-02,1.696479879319667816e-02,4.061945155262947083e-02,9.832332842051982880e-03,-3.694023191928863525e-02,-7.249249611049890518e-03,3.261747956275939941e-01,8.921848982572555542e-02,8.062155544757843018e-02,-3.506596386432647705e-02,-6.010903790593147278e-02,2.321888059377670288e-01,5.043131485581398010e-02,1.600989326834678650e-02,-1.147106289863586426e-01,8.907088637351989746e-02,-1.866739094257354736e-01,-1.688175201416015625e-01,-2.710479795932769775e-01,-1.594576239585876465e-02,-2.542634010314941406e-01,-2.836327068507671356e-02,-3.412316739559173584e-02,-1.255498975515365601e-01,-1.390765160322189331e-01,1.710339188575744629e-01,2.093050926923751831e-01,6.095051169395446777e-01,1.374952942132949829e-01,-4.103749394416809082e-01,-7.998330593109130859e-01,-6.863150000572204590e-01,-2.273800969123840332e-01,3.125610947608947754e-01,9.971548616886138916e-02,2.544522983953356743e-03,5.460501834750175476e-02,1.828952282667160034e-01,2.475388348102569580e-01,4.008584618568420410e-01,4.839259684085845947e-01,2.970970571041107178e-01,5.186368897557258606e-02,-2.399893105030059814e-02,-1.051887124776840210e-02,1.996577233076095581e-01,-6.834598723798990250e-03,-2.528696656227111816e-01,4.676536470651626587e-02,-2.436676174402236938e-01,1.277399957180023193e-01,-6.713785976171493530e-02,-1.005278676748275757e-01,1.584491580724716187e-01,-1.234629824757575989e-01,8.769094944000244141e-02,3.416405990719795227e-02,-4.283208772540092468e-02,2.344871908426284790e-01,1.014486178755760193e-01,1.401782184839248657e-01,2.146488428115844727e-01,1.304198428988456726e-02,6.002254318445920944e-03,2.170141190290451050e-01,1.675467006862163544e-02,6.632111966609954834e-02,8.814103901386260986e-02,1.642162352800369263e-01,4.872024804353713989e-02,6.645156443119049072e-02,7.112774252891540527e-02,-1.758487969636917114e-01,-1.276724226772785187e-02,-2.332994788885116577e-01,-1.236949935555458069e-01,-5.335295200347900391e-02,-2.259743213653564453e-02,-8.936194330453872681e-02,-1.996752619743347168e-01,-2.980409860610961914e-01,1.298292279243469238e-01,-1.961565911769866943e-01,-1.373527646064758301e-01,-1.170062497258186340e-01,2.007386274635791779e-02,-2.223681658506393433e-01,1.088190153241157532e-01,-8.935938030481338501e-02,1.998950392007827759e-01,-2.371882647275924683e-01,1.240669339895248413e-01,2.102467566728591919e-01,3.502171114087104797e-02,1.444858033210039139e-02,-3.670458868145942688e-02,-1.959129236638545990e-02,-5.229377374053001404e-02,2.132512032985687256e-01,-2.706399559974670410e-01,-6.251662969589233398e-02,3.094583153724670410e-01,1.015306413173675537e-01,-1.666277050971984863e-01,1.723574399948120117e-01,1.443410385400056839e-02,1.633975096046924591e-02,1.048951074481010437e-01,-5.844052135944366455e-02,-2.103029489517211914e-01,7.141897827386856079e-02,-3.687634691596031189e-02,-8.374519646167755127e-03,-8.475607633590698242e-02,5.346982553601264954e-02,-2.925288677215576172e-02,6.818628869950771332e-03,-3.495411202311515808e-02,2.055319398641586304e-01,-5.484885722398757935e-02,-2.362223342061042786e-02,1.260798871517181396e-01,2.347565591335296631e-01,6.652942299842834473e-02,3.566818311810493469e-02,-1.815397739410400391e-01,2.656013071537017822e-01,1.442363262176513672e-01,1.107212156057357788e-01,1.245565265417098999e-01,5.845645815134048462e-02,1.101179271936416626e-01,-4.032848868519067764e-03,6.051502376794815063e-02,1.558720767498016357e-01,4.499430209398269653e-02,4.668035358190536499e-02,-4.180802777409553528e-02,1.864741891622543335e-01,2.315512597560882568e-01,-2.152080088853836060e-01,7.142728567123413086e-02,-6.659574061632156372e-02,-2.138736471533775330e-02,7.591248303651809692e-02,-1.252763271331787109e-01,-5.719149485230445862e-02,-2.375538460910320282e-02,-4.376775398850440979e-02,2.491829246282577515e-01,-7.301020435988903046e-03,3.019623756408691406e-01,1.028715819120407104e-01,1.638129502534866333e-01,4.403147995471954346e-01,3.016012310981750488e-01,4.820407927036285400e-01,8.908875584602355957e-01,1.076643228530883789e+00,1.034121632575988770e+00,3.484280109405517578e-01,-2.828698754310607910e-01,1.374314278364181519e-01,-1.395027637481689453e-01,-1.374910399317741394e-02,9.238874167203903198e-02,-2.135160267353057861e-01,-4.701025784015655518e-01,-1.236748397350311279e-01,-5.804568901658058167e-02,2.037856727838516235e-01,6.526204943656921387e-02,2.147448211908340454e-01,-1.643889956176280975e-02,1.533479541540145874e-01,-2.879021465778350830e-01,3.020270168781280518e-01,1.116662099957466125e-02,1.682289540767669678e-01,4.479067027568817139e-02,1.601830422878265381e-01,3.718507289886474609e-02,2.100753039121627808e-01,9.678202122449874878e-02,-6.307165324687957764e-02,1.153347343206405640e-01,-1.343383789062500000e-01,4.986038058996200562e-02,2.430895715951919556e-02,2.326525896787643433e-01,-1.682841777801513672e-02,3.865123391151428223e-01,1.714941263198852539e-01,1.273024529218673706e-01,4.226272106170654297e-01,5.901820585131645203e-02,2.157202735543251038e-02,1.394862681627273560e-01,1.708474904298782349e-01,-3.144137561321258545e-02,-1.176775842905044556e-01,1.949597150087356567e-01,1.235100701451301575e-01,6.101825088262557983e-02,2.823488414287567139e-01,-6.723839044570922852e-02,1.994588375091552734e-01,-3.613048419356346130e-02,1.248180642724037170e-01,1.227694302797317505e-01,-6.321420520544052124e-02,-2.292032390832901001e-01,2.677085101604461670e-01,-2.080726921558380127e-01,1.516375988721847534e-01,-3.273799121379852295e-01,-8.894583582878112793e-02,-3.623256459832191467e-03,-8.429124951362609863e-02,-2.883797883987426758e-02,9.620042145252227783e-02,1.110076624900102615e-02,1.663226634263992310e-01,-3.266633152961730957e-01,1.593310385942459106e-01,-9.437380731105804443e-02,8.161070197820663452e-02,-2.736565470695495605e-01,2.878732681274414062e-01,-1.112117916345596313e-01,-9.875625371932983398e-02,-1.156418677419424057e-02,9.063020348548889160e-02,2.561284899711608887e-01,-3.108299970626831055e-01,-2.707345597445964813e-02,-3.934164345264434814e-02,1.053491681814193726e-01,8.205415308475494385e-02,-4.058752581477165222e-02,8.152247965335845947e-02,-3.726951032876968384e-02,-1.444208621978759766e-01,-1.479312926530838013e-01,-7.097167521715164185e-02,6.677260994911193848e-02,-2.081320285797119141e-01,1.173385083675384521e-01,-2.340622842311859131e-01,-8.271913975477218628e-02,-8.936296403408050537e-02,-2.774050533771514893e-01,-1.410001218318939209e-01,-2.653214931488037109e-01,-8.686247467994689941e-02,2.409259416162967682e-02,5.987335462123155594e-03,-2.969050705432891846e-01,-3.003840148448944092e-01,-4.027287289500236511e-02,-2.436672449111938477e-01,-1.416626721620559692e-01,-1.057720929384231567e-01,-1.804069280624389648e-01,-3.560366854071617126e-02,2.523477887734770775e-03,-1.808304935693740845e-01,5.344371497631072998e-02,-1.285259872674942017e-01,-1.476604491472244263e-03,3.813998773694038391e-02,-9.371304512023925781e-02,-1.905046254396438599e-01,-1.188737303018569946e-01,-2.030851840972900391e-01,-2.089905291795730591e-01,-3.478674590587615967e-02,2.427276223897933960e-02,-9.043691307306289673e-02,-8.503885939717292786e-03,1.044799387454986572e-01,4.606474936008453369e-02,6.688322406262159348e-03,3.000209629535675049e-01,3.477095812559127808e-02,-4.720489084720611572e-01,-1.889443844556808472e-01,-6.301125288009643555e-01,3.710375726222991943e-01,1.356829404830932617e-01,-5.437510609626770020e-01,4.242736473679542542e-02,1.764951460063457489e-02,-9.155006706714630127e-02,1.532782316207885742e-01,4.455626010894775391e-01,1.254330128431320190e-01,-6.475642919540405273e-01,-2.332893345737829804e-04,4.564627632498741150e-02,6.004521623253822327e-03,-1.167694777250289917e-01,1.821722388267517090e-01,-1.230958774685859680e-01,1.754658296704292297e-02,2.484394237399101257e-02,-1.834124512970447540e-02,-5.750441551208496094e-02,1.023773699998855591e-01,-1.591761261224746704e-01,-1.756418794393539429e-01,1.814141571521759033e-01,-2.531743347644805908e-01,1.087348610162734985e-01,1.823647320270538330e-02,1.259198784828186035e-01,-1.145301461219787598e-01,1.570597290992736816e-01,5.685625365003943443e-04,6.317440420389175415e-02,3.076305054128170013e-02,-5.021958798170089722e-02,-1.062293071299791336e-02,-1.036369204521179199e-01,-9.724067896604537964e-02,-1.414496749639511108e-01,-1.730241328477859497e-01,5.060108006000518799e-02,-2.642138600349426270e-01,1.112188547849655151e-01,-2.775413356721401215e-02,-2.674070298671722412e-01,2.736236900091171265e-02,-9.639108926057815552e-02,-6.309455633163452148e-02,-5.791650712490081787e-02,4.861479252576828003e-02,-3.893588483333587646e-01,1.154051348567008972e-01,1.219317466020584106e-01,-2.334832586348056793e-02,-2.486397325992584229e-02,9.096187353134155273e-02,-2.868581376969814301e-02,-7.355881482362747192e-02,-5.300847813487052917e-02,1.691522002220153809e-01,1.468248963356018066e-01,1.610121577978134155e-01,2.833892777562141418e-02,4.048402607440948486e-02,-1.642517372965812683e-02,-4.709597304463386536e-02,-4.173983633518218994e-02,7.075409591197967529e-02,-2.305503487586975098e-01,8.670388907194137573e-02,-6.608489900827407837e-02,-1.143736988306045532e-01,2.249791622161865234e-01,-1.875443905591964722e-01,9.636589884757995605e-02,1.492943763732910156e-01,-1.685556210577487946e-02,1.500148028135299683e-01,-4.795838892459869385e-02,1.266682520508766174e-03,-2.104107439517974854e-01,2.305121570825576782e-01,-3.906864300370216370e-02,8.325619995594024658e-02,5.161553993821144104e-02,-2.565397508442401886e-02,7.323236763477325439e-02,-2.124835103750228882e-01,1.262219846248626709e-01,8.283510804176330566e-02,-2.020523510873317719e-02,3.951523825526237488e-02,-1.961410343647003174e-01,-4.655599594116210938e-03,2.320713922381401062e-02,1.138198226690292358e-01,5.377323552966117859e-02,-1.632544212043285370e-02,1.719584912061691284e-01,1.747659966349601746e-02,7.810550928115844727e-02,8.450243622064590454e-02,-2.209635078907012939e-02,2.567875683307647705e-01,6.742402166128158569e-02,4.958034679293632507e-02,7.317169755697250366e-02,1.440111249685287476e-01,8.749886415898799896e-03,7.327260822057723999e-02,5.494336411356925964e-02,1.762660741806030273e-01,-3.393714129924774170e-01,1.031218469142913818e-01,2.988953329622745514e-02,-2.885070741176605225e-01,1.351652592420578003e-01,-1.832389980554580688e-01,4.474182426929473877e-02,-1.047549992799758911e-01,1.771310120820999146e-01,-5.318999662995338440e-02,1.702992320060729980e-01,1.061265990138053894e-01,-2.057017683982849121e-01,9.157256782054901123e-02,9.775456190109252930e-01,-5.020269155502319336e-01,-1.213995575904846191e+00,-1.922353208065032959e-01,6.432948708534240723e-01,-1.628638952970504761e-01,1.873723417520523071e-01,5.189436301589012146e-02,-4.370671510696411133e-02,2.086433023214340210e-02,1.063976213335990906e-01,3.996263146400451660e-01,5.805407762527465820e-01,6.598107814788818359e-01,3.068324625492095947e-01,-1.899924278259277344e-01,-3.640911579132080078e-01,-1.804623603820800781e-01,-2.087770849466323853e-01,2.626442611217498779e-01,7.685555610805749893e-03,8.876366168260574341e-02,1.110745295882225037e-01,1.116781532764434814e-01,6.142556667327880859e-02,2.980217039585113525e-01,-1.641275584697723389e-01,-7.261955738067626953e-02,-1.121509447693824768e-01,2.915466763079166412e-02,-1.244988292455673218e-01,1.179000735282897949e-01,1.039562895894050598e-01,-1.522551383823156357e-02,1.729858368635177612e-01,-9.479548782110214233e-02,1.022709384560585022e-01,1.962574422359466553e-01,-1.521902084350585938e-01,-1.025559976696968079e-01,1.703269034624099731e-02,-2.228298485279083252e-01,-1.511410623788833618e-01,-4.496345669031143188e-02,2.457413375377655029e-01,-2.421398647129535675e-02,-6.045798584818840027e-02,1.481286436319351196e-01,-1.282488554716110229e-01,2.356279045343399048e-01,-1.895170658826828003e-01,6.646373122930526733e-02,3.374538570642471313e-02,2.143300324678421021e-01,-2.618934400379657745e-02,-4.783385619521141052e-02,-6.593087315559387207e-02,1.694520562887191772e-01,-3.525966778397560120e-02,-2.124544829130172729e-01,-1.530319899320602417e-01,-8.294271305203437805e-03,-1.367495208978652954e-01,1.313542872667312622e-01,-1.544182151556015015e-01,2.210290543735027313e-02,-1.512364298105239868e-01,1.640799641609191895e-02,-1.302477717399597168e-01,-3.234290778636932373e-01,1.751894876360893250e-02,-1.783155836164951324e-02,-2.917457818984985352e-01,1.333675980567932129e-01,-2.205967158079147339e-01,-2.379610687494277954e-01,-2.640574574470520020e-01,-1.594085097312927246e-01,-1.995062679052352905e-01,-4.005570411682128906e-01,-2.748273126780986786e-02,-1.659376472234725952e-01,-5.694710090756416321e-02,-1.880350857973098755e-01,2.186899483203887939e-01,-3.549894690513610840e-01,-7.079555839300155640e-02,-1.275358200073242188e-01,1.574794948101043701e-01,-2.803672477602958679e-02,-2.377145737409591675e-01,1.362416706979274750e-02,-1.986001729965209961e-01,-1.815643161535263062e-02,-1.209023408591747284e-03,-1.320183426141738892e-01,-1.383758783340454102e-01,-9.777268767356872559e-02,-1.909340918064117432e-02,-5.221679806709289551e-01,-1.125404015183448792e-01,-1.177368834614753723e-01,1.297007352113723755e-01,-1.301951706409454346e-01,-1.278174966573715210e-01,1.047630161046981812e-01,-4.455406367778778076e-01,-3.832527101039886475e-01,-6.748855113983154297e-02,-1.166951954364776611e-01,5.291669070720672607e-02,-1.539249420166015625e-01,-1.632364690303802490e-01,-2.165318280458450317e-02,-2.156953811645507812e-01,-2.239940315485000610e-01,-1.234560087323188782e-01,-8.787037432193756104e-02,-5.122143030166625977e-02,-2.155595272779464722e-01,-3.857845366001129150e-01,-1.679582893848419189e-01,-1.931173652410507202e-01,-8.917932212352752686e-02,-3.869064748287200928e-01,-5.070832371711730957e-01,-7.162033319473266602e-01,-2.092117443680763245e-02,5.817858576774597168e-01,8.626950979232788086e-01,3.773127198219299316e-01,2.199253588914871216e-01,-9.600409120321273804e-02,-2.924684286117553711e-01,7.960630953311920166e-02,1.803437992930412292e-02,4.013359248638153076e-01,6.578344851732254028e-02,4.677884578704833984e-01,5.084300041198730469e-01,6.589195132255554199e-01,5.645632743835449219e-01,-9.033846110105514526e-02,-1.023473739624023438e-01,-2.641594111919403076e-01,-1.967756748199462891e-01,2.665390074253082275e-02,4.174790531396865845e-02,-7.341135293245315552e-02,3.594217821955680847e-02,1.749960482120513916e-01,-1.386985629796981812e-01,-5.337475985288619995e-02,1.670285910367965698e-01,1.864401400089263916e-01,6.378769129514694214e-02,1.721713244915008545e-01,2.401428818702697754e-01,-1.050892751663923264e-05,2.215677499771118164e-01,3.193785548210144043e-01,1.159472092986106873e-01,1.922091841697692871e-01,2.770194113254547119e-01,1.937408298254013062e-01,4.129390418529510498e-02,3.310315012931823730e-01,4.900243505835533142e-02,3.291935101151466370e-02,2.480874806642532349e-01,-5.890173465013504028e-02,4.375592470169067383e-01,7.739770412445068359e-02,-1.995202153921127319e-01,2.134999930858612061e-01,4.329457879066467285e-02,1.986420750617980957e-01,2.087445855140686035e-01,5.266129598021507263e-02,9.829191118478775024e-02,6.310434639453887939e-02,9.373777359724044800e-02,2.004285752773284912e-01,-1.803617551922798157e-02,2.751266956329345703e-01,-8.903688192367553711e-02,8.714333921670913696e-02,-2.983630076050758362e-02,-9.099337458610534668e-02,2.162892371416091919e-01,-1.631713509559631348e-01,1.815034598112106323e-01,2.805472016334533691e-01,1.418591588735580444e-01,2.538378536701202393e-01,1.145971044898033142e-01,3.486383706331253052e-03,-2.155823458451777697e-04,2.273340225219726562e-01,-8.160571008920669556e-02,2.199229896068572998e-01,-4.545003920793533325e-02,1.695907264947891235e-01,6.749056279659271240e-02,-1.859041489660739899e-02,1.039044931530952454e-01,9.164246730506420135e-03,1.200607568025588989e-01,1.971387565135955811e-01,3.395849764347076416e-01,3.441621363162994385e-01,-9.719005972146987915e-02,-9.331077337265014648e-02,-2.365237772464752197e-01,6.753495335578918457e-02,-1.168387010693550110e-01,8.741349726915359497e-02,2.665361389517784119e-03,2.302631586790084839e-01,2.086380571126937866e-01,1.610052436590194702e-01,-8.872558176517486572e-02,2.714837715029716492e-02,1.136632263660430908e-01,1.339196413755416870e-01,4.859771952033042908e-02,-1.901242285966873169e-01,-1.817880943417549133e-02,7.116610556840896606e-02,4.787271097302436829e-02,2.780577838420867920e-01,1.662866175174713135e-01,-6.559637933969497681e-02,2.091466635465621948e-01,2.381326556205749512e-01,2.397965341806411743e-01,4.253844618797302246e-01,3.474072217941284180e-01,5.688328528776764870e-04,2.988641262054443359e-01,3.813372924923896790e-02,3.260830938816070557e-01,3.259825110435485840e-01,3.252751529216766357e-01,7.606568187475204468e-02,2.795296609401702881e-01,2.792639434337615967e-01,3.567915856838226318e-01,-1.119957044720649719e-01,3.141587376594543457e-01,2.390747815370559692e-01,-1.142132133245468140e-01,-1.351258158683776855e-01,7.373269647359848022e-02,-1.843410730361938477e-02,-1.133186370134353638e-01,-9.776608943939208984e-01,-6.960154771804809570e-01,-1.710878908634185791e-01,5.772772431373596191e-01,5.887348055839538574e-01,2.149498164653778076e-01,-2.465178258717060089e-02,9.382885694503784180e-02,2.579117380082607269e-02,-1.533512305468320847e-02,-1.968014091253280640e-01,-4.476780295372009277e-01,-3.894922137260437012e-01,-9.807427972555160522e-02,-1.542986184358596802e-01,8.626941591501235962e-02,-2.130418717861175537e-01,-2.446152120828628540e-01,-2.003467082977294922e-01,-3.955094516277313232e-02,-7.331430166959762573e-02,-1.248868107795715332e-01,-1.070564314723014832e-01,7.105068862438201904e-02,-6.475935131311416626e-02,-1.794315725564956665e-01,-9.516783803701400757e-02,-1.003110557794570923e-01,-1.254691034555435181e-01,-8.023717254400253296e-02,2.704606624320149422e-03,-6.364504992961883545e-02,-1.206681653857231140e-01,7.623519003391265869e-02,1.326788216829299927e-01,-7.795851677656173706e-02,2.094782441854476929e-01,-1.819966137409210205e-01,8.278376609086990356e-02,-1.488421708345413208e-01,-6.112342700362205505e-02,-1.795193403959274292e-01,7.645993679761886597e-02,-1.208675280213356018e-01,1.481667309999465942e-01,5.024204403162002563e-02,5.905196443200111389e-02,2.607189416885375977e-01,5.375811085104942322e-02,1.961511000990867615e-02,-1.585835218429565430e-02,-4.003611952066421509e-02,-1.066681221127510071e-01,8.766520768404006958e-02,1.389352232217788696e-01,6.889014691114425659e-02,-7.694721966981887817e-02,2.183835506439208984e-01,-7.202729582786560059e-02,-2.627655863761901855e-01,-9.519518166780471802e-02,3.196633234620094299e-02,-1.002400368452072144e-02,1.716046780347824097e-01,-2.596682682633399963e-02,-1.831363290548324585e-01,3.118706401437520981e-03,7.088187616318464279e-03,-7.274815440177917480e-02,-4.786931350827217102e-02,1.783335208892822266e-01,-5.127536877989768982e-02,-4.180839657783508301e-02,-8.335531502962112427e-02,2.959171682596206665e-02,-6.597356405109167099e-04,7.905938662588596344e-03,1.435800790786743164e-01,-4.981091246008872986e-02,3.145133331418037415e-02,-1.001730337738990784e-01,8.781793527305126190e-03,-2.131903171539306641e-01,5.848648143000900745e-04,1.879484802484512329e-01,-1.082822531461715698e-01,-4.615236818790435791e-02,-4.197381809353828430e-02,-2.161490265280008316e-03,-7.920632511377334595e-02,-9.892947226762771606e-02,4.736595228314399719e-02,-7.332307100296020508e-02,-1.036864332854747772e-02,-4.142526164650917053e-02,-6.426475197076797485e-02,-6.862074136734008789e-02,2.273183781653642654e-03,-2.945895195007324219e-01,-1.530423015356063843e-01,-1.032201647758483887e-01,6.150968372821807861e-02,-1.560306549072265625e-02,7.088156044483184814e-02,-1.382834464311599731e-01,8.165816776454448700e-03,1.641557086259126663e-03,-1.241371706128120422e-01,-7.477407902479171753e-02,-2.718734182417392731e-02,-1.351521611213684082e-01,3.530584275722503662e-02,-1.029962152242660522e-01,-5.603168532252311707e-02,4.330096766352653503e-02,1.206409744918346405e-02,-3.163906186819076538e-02,-4.078555107116699219e-02,-2.163390628993511200e-02,-1.740864962339401245e-01,-1.404804289340972900e-01,-1.070955768227577209e-01,-1.023654341697692871e-01,-1.100936159491539001e-01,4.699543863534927368e-02,-1.856247037649154663e-01,5.750858411192893982e-02,-3.417935669422149658e-01,-5.114267468452453613e-01,-6.354480981826782227e-01,-2.083954066038131714e-01,8.292791247367858887e-01,5.593308210372924805e-01,-1.086789742112159729e-02,4.364158213138580322e-01,2.439146786928176880e-01,8.797269314527511597e-02,-4.123153090476989746e-01,-6.411705613136291504e-01,-4.640594422817230225e-01,4.909923672676086426e-02,4.620004296302795410e-01,6.273531317710876465e-01,6.381242275238037109e-01,4.495024979114532471e-01,1.708534061908721924e-01,-8.297723531723022461e-02,2.164040803909301758e-01,-2.152917087078094482e-01,-2.344172820448875427e-02,2.677348814904689789e-02,1.673585474491119385e-01,1.863789856433868408e-01,1.426559388637542725e-01,-1.804365962743759155e-01,3.073042929172515869e-01,7.030688971281051636e-02,2.593251168727874756e-01,-6.096096336841583252e-02,1.890840679407119751e-01,1.146998107433319092e-01,-1.632943302392959595e-01,3.437643647193908691e-01,9.792937897145748138e-03,-7.311093062162399292e-02,1.097134947776794434e-01,2.834325134754180908e-01,-1.725747585296630859e-01,-1.061447784304618835e-01,2.381650209426879883e-01,1.114237681031227112e-01,4.126203432679176331e-02,2.123482823371887207e-01,1.176885366439819336e-01,-4.913858138024806976e-03,-1.104761734604835510e-01,-4.726231470704078674e-02,-1.687216758728027344e-01,2.883225381374359131e-01,7.091572135686874390e-02,-1.142567396163940430e-01,1.377005279064178467e-01,3.441967070102691650e-01,-1.097471192479133606e-01,-8.021975308656692505e-02,-8.821664378046989441e-03,9.118369780480861664e-04,-1.076869666576385498e-01,1.683827638626098633e-01,2.547218464314937592e-03,-3.095155656337738037e-01,1.128660589456558228e-01,8.543545007705688477e-02,6.571216136217117310e-02,-7.407327182590961456e-03,-4.592308998107910156e-01,1.460091173648834229e-01,2.450209110975265503e-01,-1.742016226053237915e-01,-1.161962300539016724e-01,1.720979213714599609e-01,-2.697578072547912598e-01,-2.030574083328247070e-01,1.311619281768798828e-01,-5.497367680072784424e-02,1.860131160356104374e-04,1.519380062818527222e-01,1.188764795660972595e-01,-3.253951966762542725e-01,1.732712388038635254e-01,-1.286369413137435913e-01,4.377307742834091187e-02,-3.247852623462677002e-02,-2.931863367557525635e-01,2.026992589235305786e-01,-2.057525366544723511e-01,2.468642443418502808e-01,-2.140765041112899780e-01,2.604442238807678223e-01,-8.379048854112625122e-02,2.491413056850433350e-01,2.111393772065639496e-02,-1.396833658218383789e-01,-2.941420078277587891e-01,2.223598062992095947e-01,-2.084284722805023193e-01,8.226880431175231934e-02,-3.425249829888343811e-02,9.798914939165115356e-02,-1.299363374710083008e-01,-2.046712189912796021e-01,-1.279760897159576416e-01,8.526203781366348267e-02,3.470331197604537010e-03,-2.358607053756713867e-01,-3.637116774916648865e-02,-1.150849536061286926e-01,1.935552656650543213e-01,-2.515639737248420715e-02,-1.132180020213127136e-01,1.277035027742385864e-01,3.153889253735542297e-02,-2.150217592716217041e-01,4.269119352102279663e-02,-2.948800325393676758e-01,1.146650612354278564e-01,-1.045946106314659119e-01,1.713913977146148682e-01,-6.776275485754013062e-02,-2.541815638542175293e-01,-2.284491658210754395e-01,1.703607104718685150e-02,1.735707521438598633e-01,1.033389195799827576e-01,4.513218104839324951e-01,8.744094520807266235e-02,-4.277203679084777832e-01,-3.323228657245635986e-01,-2.111718505620956421e-01,7.421076297760009766e-02,-3.363586589694023132e-02,-2.225661873817443848e-01);
    constant w1r_imag : w1r_array := (1.048476099967956543e-01,-8.256702870130538940e-02,2.556248307228088379e-01,1.123163700103759766e+00,3.380401730537414551e-01,-1.075198888778686523e+00,-3.591450750827789307e-01,5.709412097930908203e-01,2.626438438892364502e-01,1.141354888677597046e-01,3.031064383685588837e-02,3.484052047133445740e-02,-1.179515495896339417e-01,-5.397621914744377136e-02,-1.568792909383773804e-01,-1.362563222646713257e-01,-1.008177623152732849e-01,-9.887901693582534790e-02,1.054204702377319336e-01,-2.071048170328140259e-01,5.881117284297943115e-02,2.800940722227096558e-02,-4.979359731078147888e-02,-2.043791860342025757e-01,2.589261233806610107e-01,-7.725502550601959229e-02,-1.828214973211288452e-01,-6.599551439285278320e-02,-2.070333361625671387e-01,-6.313651800155639648e-02,-1.184800788760185242e-01,8.541505038738250732e-02,-2.058770060539245605e-01,1.103430762887001038e-01,-5.669205449521541595e-03,8.737081289291381836e-02,1.624223887920379639e-01,-1.330325454473495483e-01,6.737295538187026978e-02,-5.988926067948341370e-02,4.832535982131958008e-02,-2.462885528802871704e-02,-2.653828561305999756e-01,2.140373736619949341e-01,-3.004642724990844727e-01,-1.425092071294784546e-01,-1.413750648498535156e-01,2.170896157622337341e-02,-1.747413724660873413e-01,4.333593323826789856e-02,-6.055524200201034546e-02,-2.490895390510559082e-01,-3.877251595258712769e-02,-3.779453337192535400e-01,5.749313859269022942e-04,-1.859906762838363647e-01,2.204531133174896240e-01,7.211564481258392334e-02,-1.071118116378784180e-01,-6.679744273424148560e-02,-3.069089492782950401e-03,5.411431938409805298e-02,9.909652173519134521e-02,-4.132999107241630554e-02,3.289183229207992554e-02,2.696004882454872131e-02,2.611870411783456802e-03,-2.275773286819458008e-01,-1.175285652279853821e-01,-1.635852269828319550e-02,-3.445752561092376709e-01,-3.126559033989906311e-02,-3.088084980845451355e-03,2.202566415071487427e-01,-5.239449739456176758e-01,-1.454411260783672333e-02,-1.979403048753738403e-01,2.179197669029235840e-01,-2.115653008222579956e-01,-1.460226774215698242e-01,-2.760922610759735107e-01,-3.192843198776245117e-01,8.821115642786026001e-02,-1.335728168487548828e-02,-1.653667539358139038e-01,-1.008450910449028015e-01,1.934038400650024414e-01,-3.115113941021263599e-04,1.877135187387466431e-01,1.856458783149719238e-01,4.264616966247558594e-02,3.462217003107070923e-02,6.063042208552360535e-03,-7.357682287693023682e-02,1.455942690372467041e-01,2.048266306519508362e-02,-1.558424532413482666e-01,1.027707532048225403e-01,7.106177508831024170e-02,3.194089606404304504e-02,3.451138362288475037e-02,4.668652266263961792e-02,2.213485352694988251e-02,2.306721061468124390e-01,6.642984598875045776e-02,4.165827631950378418e-01,4.412837792187929153e-03,4.991354420781135559e-02,1.180797889828681946e-01,3.118959963321685791e-01,-1.016847118735313416e-01,2.524049580097198486e-01,-5.112317577004432678e-02,-5.125372484326362610e-02,-7.645468413829803467e-02,5.026660487055778503e-02,1.591715514659881592e-01,1.904671639204025269e-01,3.300070017576217651e-02,2.842067182064056396e-01,-1.404473483562469482e-01,4.493639469146728516e-01,1.663897484540939331e-01,-3.444250226020812988e-01,-2.968108952045440674e-01,2.638439834117889404e-01,-1.456619203090667725e-01,3.533281683921813965e-01,7.681042701005935669e-02,1.099402606487274170e-01,-6.166373938322067261e-02,1.272893995046615601e-01,4.701813682913780212e-02,3.736961185932159424e-01,-4.732147604227066040e-02,-2.966217696666717529e-02,-1.600564569234848022e-01,-2.159224264323711395e-02,-9.446694515645503998e-03,2.379530519247055054e-01,-1.004985794425010681e-01,1.162935718894004822e-01,8.812091499567031860e-02,-4.849289357662200928e-02,7.322502881288528442e-02,-7.872461341321468353e-03,1.806951314210891724e-01,-9.118878096342086792e-02,1.358621865510940552e-01,1.794659197330474854e-01,2.155326120555400848e-02,1.138077303767204285e-01,1.435897648334503174e-01,-1.664462685585021973e-02,4.356233403086662292e-02,-1.772158443927764893e-01,-1.125398129224777222e-01,1.851005703210830688e-01,-3.752737864851951599e-02,1.079671308398246765e-01,1.064243074506521225e-02,1.204488873481750488e-01,-4.468765109777450562e-02,-1.207368820905685425e-01,5.479053780436515808e-02,-1.409086436033248901e-01,-3.776707872748374939e-02,-4.583669453859329224e-02,-1.042278558015823364e-01,1.837974227964878082e-02,-1.207710951566696167e-01,-1.700441688299179077e-01,-2.426107525825500488e-01,-1.306776553392410278e-01,-1.966302394866943359e-01,5.513650551438331604e-02,-4.592053592205047607e-02,2.042176574468612671e-02,-4.899121448397636414e-02,2.268486656248569489e-02,-1.641243398189544678e-01,7.223081588745117188e-02,2.188016772270202637e-01,1.426058262586593628e-01,-6.793908774852752686e-02,5.784250795841217041e-02,-1.951034180819988251e-02,9.952615946531295776e-02,-2.552263736724853516e-01,1.239707693457603455e-02,-2.033086493611335754e-02,6.176085025072097778e-02,7.647546380758285522e-02,1.203275844454765320e-01,4.522482678294181824e-02,2.102124504745006561e-02,9.494892507791519165e-02,9.644559770822525024e-02,-6.961961276829242706e-03,8.997984230518341064e-03,1.117987483739852905e-01,2.311787605285644531e-01,-1.739659011363983154e-01,-8.307666517794132233e-03,-4.510214924812316895e-02,2.243200838565826416e-01,1.265579313039779663e-01,2.392418682575225830e-01,-1.360403895378112793e-01,2.737720608711242676e-01,2.328425273299217224e-02,3.045643568038940430e-01,5.922083184123039246e-02,3.223962187767028809e-01,-3.398337634280323982e-03,1.811007559299468994e-01,1.388596147298812866e-01,8.572813868522644043e-02,3.020089119672775269e-02,7.101635634899139404e-02,1.942358314990997314e-01,1.262495815753936768e-01,1.748176664113998413e-01,7.355145364999771118e-02,-9.830266935750842094e-04,1.949922591447830200e-01,1.728544384241104126e-01,2.335757911205291748e-01,6.190476939082145691e-02,1.496393382549285889e-01,1.649865210056304932e-01,-1.168797984719276428e-01,1.293866634368896484e-01,8.953868597745895386e-02,1.123237386345863342e-01,5.738677084445953369e-02,1.011078506708145142e-01,-1.334509160369634628e-02,2.042151689529418945e-01,8.103328943252563477e-02,3.703827038407325745e-02,-2.737531960010528564e-01,3.139300048351287842e-01,6.638650596141815186e-02,-1.680859029293060303e-01,3.456231653690338135e-01,1.181004792451858521e-01,1.845659464597702026e-01,-1.708428263664245605e-01,2.451441884040832520e-01,1.253477782011032104e-01,1.148881092667579651e-01,-1.932566910982131958e-01,-7.637030631303787231e-02,4.506660699844360352e-01,-4.307482242584228516e-01,-2.525469660758972168e-01,6.157757341861724854e-02,8.572485297918319702e-02,5.277867913246154785e-01,-4.990996122360229492e-01,-4.580484032630920410e-01,2.566319704055786133e-01,-2.378209978342056274e-01,1.030654609203338623e-01,1.071327105164527893e-01,1.188064217567443848e-01,-7.127065956592559814e-02,-6.245645694434642792e-03,-6.862635165452957153e-02,-8.129227906465530396e-02,4.731093347072601318e-02,-2.149491012096405029e-02,4.311650525778532028e-03,1.746195554733276367e-01,-7.189323753118515015e-02,-2.109613269567489624e-02,7.818286865949630737e-02,-4.675434157252311707e-02,1.854055002331733704e-02,-6.134924292564392090e-02,-1.899001002311706543e-01,-2.790644206106662750e-02,5.674408003687858582e-02,-4.214000701904296875e-02,-4.464111104607582092e-02,8.554530143737792969e-02,7.314392924308776855e-02,-1.273091137409210205e-01,-1.195553410798311234e-02,1.316679120063781738e-01,-3.629919141530990601e-02,3.358035534620285034e-02,-1.524699386209249496e-02,1.370912790298461914e-01,-1.305137425661087036e-01,-1.072886958718299866e-01,4.771887138485908508e-02,1.429355517029762268e-02,-1.897265464067459106e-01,6.319156847894191742e-03,-8.313591778278350830e-02,6.776269874535501003e-04,2.039013057947158813e-01,1.815403252840042114e-02,-5.872511491179466248e-02,1.175573319196701050e-01,-9.436856210231781006e-02,1.088828295469284058e-01,2.069654017686843872e-01,5.181772634387016296e-02,1.935623437166213989e-01,3.301637768745422363e-01,9.973010420799255371e-02,-7.607162930071353912e-03,-2.872395142912864685e-02,1.499052252620458603e-02,-9.293343126773834229e-02,-2.522112131118774414e-01,2.363964766263961792e-01,2.594094574451446533e-01,1.060309484601020813e-01,1.995236426591873169e-02,3.157444894313812256e-01,4.367461428046226501e-02,-7.125858962535858154e-02,-3.781617060303688049e-02,-1.263412181288003922e-02,1.163768116384744644e-02,-3.812214732170104980e-02,-6.996574997901916504e-02,2.794980108737945557e-01,-6.960454583168029785e-02,-3.472932428121566772e-02,2.972398400306701660e-01,4.203954711556434631e-02,5.130625888705253601e-02,-4.556823521852493286e-02,-3.341605514287948608e-02,2.529923319816589355e-01,-5.569344013929367065e-02,-5.785269290208816528e-02,7.582182437181472778e-02,-4.055120050907135010e-02,6.187034025788307190e-02,1.478412896394729614e-01,2.905069887638092041e-01,-1.074452474713325500e-01,2.835520170629024506e-02,5.350799486041069031e-02,-2.647154498845338821e-03,-2.001721970736980438e-02,-1.218446902930736542e-02,-1.257880032062530518e-01,8.824668079614639282e-02,-1.351726502180099487e-01,1.495306491851806641e-01,-1.899365931749343872e-01,1.108492910861968994e-01,-3.186919167637825012e-02,7.502502948045730591e-02,2.727946043014526367e-01,-6.452911347150802612e-02,1.336039043962955475e-02,-2.428094148635864258e-01,2.390271611511707306e-02,7.279122620820999146e-02,5.486505851149559021e-02,3.143156766891479492e-01,-7.086377590894699097e-02,9.475449472665786743e-02,2.833034694194793701e-01,1.557794027030467987e-02,-1.582555659115314484e-02,1.855603903532028198e-01,-1.128132864832878113e-01,-5.348108410835266113e-01,-2.224464714527130127e-01,-3.882160410284996033e-02,3.447489738464355469e-01,3.585999310016632080e-01,-5.550867915153503418e-01,6.793146729469299316e-01,6.780138704925775528e-03,1.551132351160049438e-01,4.464692771434783936e-01,2.395292818546295166e-01,-1.589437574148178101e-01,3.112961947917938232e-01,9.927305579185485840e-02,-6.171337515115737915e-02,9.354875981807708740e-02,-9.859264642000198364e-02,-3.073392994701862335e-02,-1.203660890460014343e-01,1.610904186964035034e-01,7.959930226206779480e-03,-1.857713758945465088e-01,1.904251128435134888e-01,9.027902781963348389e-02,1.395144760608673096e-01,-1.149459555745124817e-02,5.919200554490089417e-02,-2.812573313713073730e-01,6.075624749064445496e-02,2.234238684177398682e-01,-5.203613638877868652e-02,1.457101106643676758e-01,1.143207657150924206e-03,2.186880260705947876e-01,4.204227030277252197e-02,1.095707714557647705e-01,-5.355275049805641174e-02,2.099704146385192871e-01,-1.217155531048774719e-01,1.563641279935836792e-01,5.715837329626083374e-02,1.363315880298614502e-01,-2.083259820938110352e-01,1.793965101242065430e-01,1.968529224395751953e-01,-1.555668711662292480e-01,2.641545236110687256e-01,-1.338125616312026978e-01,-3.399381786584854126e-02,3.702575862407684326e-01,-2.554350793361663818e-01,-4.125460982322692871e-02,-1.392528712749481201e-01,-2.527339383959770203e-02,-5.944805592298507690e-02,-2.320809289813041687e-02,1.717018485069274902e-01,-1.028770431876182556e-01,5.836256965994834900e-02,-1.695198714733123779e-01,-6.914105266332626343e-02,-2.307744771242141724e-01,-7.414009422063827515e-02,6.168485805392265320e-02,-1.437803208827972412e-01,-1.031916886568069458e-01,1.000000536441802979e-01,-1.441066265106201172e-01,7.990419864654541016e-03,-2.022310644388198853e-01,-3.216045796871185303e-01,8.707571029663085938e-02,2.188525646924972534e-01,-3.442552387714385986e-01,-2.333721667528152466e-01,1.860362142324447632e-01,-6.154824793338775635e-02,-2.654877901077270508e-01,4.764740914106369019e-02,-3.024793863296508789e-01,2.015208154916763306e-01,1.657106280326843262e-01,-8.284711837768554688e-02,-1.552367061376571655e-01,-5.888041853904724121e-02,-9.104768931865692139e-02,-1.655066013336181641e-01,-4.955251142382621765e-02,-6.807813793420791626e-02,-1.374121308326721191e-01,-2.307793051004409790e-01,-1.159815639257431030e-01,9.119215607643127441e-02,-2.151127010583877563e-01,-6.512360274791717529e-02,2.093658149242401123e-01,-2.157385647296905518e-01,1.203827261924743652e-01,2.531490921974182129e-01,-1.623463332653045654e-01,2.261524349451065063e-01,6.292125582695007324e-02,4.104775190353393555e-02,3.183397352695465088e-01,7.021858543157577515e-02,1.023975387215614319e-01,1.296762675046920776e-01,2.978441119194030762e-01,1.757643222808837891e-01,6.883801519870758057e-02,2.795023322105407715e-01,7.999080419540405273e-02,-4.265860468149185181e-02,2.397063374519348145e-01,1.611277312040328979e-01,1.406133323907852173e-01,2.324845828115940094e-02,1.277594566345214844e-01,1.900013536214828491e-01,1.664846837520599365e-01,-2.149989269673824310e-02,6.401488184928894043e-02,-2.576290071010589600e-01,3.002951443195343018e-01,4.267917945981025696e-02,6.249931454658508301e-02,1.221747472882270813e-01,-1.103624552488327026e-01,-6.032945960760116577e-02,-2.024321854114532471e-01,-3.312014937400817871e-01,-4.369681477546691895e-01,-1.599870920181274414e-01,2.559682726860046387e-01,4.888711273670196533e-01,2.378984540700912476e-01,5.759409070014953613e-02,1.591315120458602905e-01,3.364555537700653076e-01,2.635127305984497070e-01,-6.581446528434753418e-01,8.315657824277877808e-02,1.867289543151855469e-01,-3.849102854728698730e-01,2.471446692943572998e-01,6.607511639595031738e-01,9.097727388143539429e-02,-4.075576737523078918e-02,2.580286264419555664e-01,-4.484649375081062317e-02,4.942898079752922058e-02,4.269012250006198883e-03,-6.800766568630933762e-03,4.737421125173568726e-02,1.571195572614669800e-02,4.072995483875274658e-02,1.188786104321479797e-01,6.874603033065795898e-02,1.820650398731231689e-01,-6.077773496508598328e-02,4.265925660729408264e-02,1.968323886394500732e-01,-4.907366260886192322e-02,9.169491380453109741e-02,-9.157065302133560181e-02,2.553522773087024689e-02,1.865414977073669434e-01,-9.288322180509567261e-02,1.269591301679611206e-01,-3.902490064501762390e-02,1.433674991130828857e-01,8.516109734773635864e-02,-5.560371279716491699e-02,2.603102289140224457e-02,5.495151504874229431e-02,7.023803144693374634e-02,-9.396569430828094482e-02,5.693755671381950378e-02,2.300235070288181305e-02,-2.283285409212112427e-01,1.795768737792968750e-01,-1.780250817537307739e-01,-6.984028499573469162e-03,-2.765939198434352875e-02,-4.453689604997634888e-02,-6.095991283655166626e-02,2.901270985603332520e-01,-1.583061814308166504e-01,-2.277905866503715515e-02,1.247892901301383972e-01,-3.159662336111068726e-02,-9.336293488740921021e-02,5.685725063085556030e-02,-1.551585495471954346e-01,1.273438241332769394e-02,-7.655496895313262939e-02,4.003074020147323608e-02,1.232973784208297729e-01,-2.514385581016540527e-01,4.429817199707031250e-02,-1.038567498326301575e-01,-1.328114569187164307e-01,-1.334230899810791016e-01,1.500649899244308472e-01,-3.447496592998504639e-01,8.838011883199214935e-03,-3.007248044013977051e-01,-2.933690845966339111e-01,8.752314001321792603e-02,3.970361500978469849e-02,-1.220484822988510132e-01,4.397930577397346497e-02,-2.090407460927963257e-01,8.676001429557800293e-02,1.050565242767333984e-01,-1.287483870983123779e-01,1.335307583212852478e-02,1.109717637300491333e-01,-1.009510383009910583e-01,2.599609270691871643e-02,-3.645411133766174316e-02,-4.820497706532478333e-02,1.696608401834964752e-02,1.090344190597534180e-01,7.136293500661849976e-02,-2.786469645798206329e-03,9.412924759089946747e-03,-8.035549521446228027e-02,1.696565002202987671e-01,2.387066334486007690e-01,2.299169898033142090e-01,1.950147561728954315e-02,3.115254640579223633e-01,4.230865836143493652e-02,1.317175626754760742e-01,6.310810148715972900e-02,7.329732924699783325e-02,5.196833983063697815e-02,-4.082811996340751648e-02,6.685417890548706055e-02,-2.360476739704608917e-02,6.897930055856704712e-03,1.113893464207649231e-01,1.858306378126144409e-01,4.237444326281547546e-02,2.238937094807624817e-02,8.009767532348632812e-02,1.266958117485046387e-01,-1.393396290950477123e-03,-2.042967379093170166e-01,5.719795357435941696e-03,-7.289048284292221069e-02,-9.375734627246856689e-02,9.423058480024337769e-02,3.440025821328163147e-02,2.571164369583129883e-01,-4.967429041862487793e-01,-5.285308957099914551e-01,1.480288505554199219e+00,1.083396553993225098e+00,-9.746512770652770996e-01,1.111074462532997131e-01,5.628814101219177246e-01,-9.041110426187515259e-02,2.334129959344863892e-01,3.869762122631072998e-01,5.068907737731933594e-01,7.394148707389831543e-01,4.479215145111083984e-01,1.398939341306686401e-01,-5.838117599487304688e-01,-4.316306710243225098e-01,-3.114469647407531738e-01,-2.347744107246398926e-01,-5.146448686718940735e-02,8.538696914911270142e-02,2.126812934875488281e-01,4.260619729757308960e-02,3.478783667087554932e-01,-2.003006935119628906e-01,7.910574204288423061e-04,-1.316177994012832642e-01,1.409418582916259766e-01,1.921612173318862915e-01,-2.195290625095367432e-01,-3.138530552387237549e-01,-1.276490837335586548e-01,3.376930356025695801e-01,-1.616248674690723419e-02,1.322513669729232788e-01,2.342125177383422852e-01,-3.948649391531944275e-03,2.195627093315124512e-01,5.930515751242637634e-02,2.718237042427062988e-01,7.163972407579421997e-02,1.941177397966384888e-01,-4.915409907698631287e-02,1.187315862625837326e-02,1.712468862533569336e-01,7.264963537454605103e-02,-2.123531252145767212e-01,5.675301421433687210e-03,2.507809549570083618e-03,-2.574164234101772308e-02,-7.165040820837020874e-02,2.033514827489852905e-01,1.311265230178833008e-01,1.337545514106750488e-01,-9.821844100952148438e-02,2.017643600702285767e-01,-1.417840421199798584e-01,2.795124053955078125e-01,-2.511397004127502441e-01,-1.216829791665077209e-01,1.283047050237655640e-01,1.455205827951431274e-01,8.396070450544357300e-02,1.249640882015228271e-01,-1.528588384389877319e-01,-2.950155921280384064e-02,2.931309640407562256e-01,-2.157266139984130859e-01,-1.602642685174942017e-01,-4.466005787253379822e-02,3.431672751903533936e-01,-1.666907519102096558e-01,6.002290546894073486e-02,2.476266622543334961e-01,-2.424401193857192993e-01,-1.901451200246810913e-01,1.273107528686523438e-01,-1.090663578361272812e-02,-9.171842038631439209e-02,-1.041674166917800903e-01,2.666364423930644989e-02,-5.239212512969970703e-01,-7.918800413608551025e-02,1.929100900888442993e-01,7.034631073474884033e-02,-4.056450352072715759e-02,2.199923433363437653e-02,-1.808238625526428223e-01,-2.311858552275225520e-04,7.812588661909103394e-02,-3.204847872257232666e-01,-6.305577605962753296e-02,1.781451851129531860e-01,-1.236917972564697266e-01,-6.889462471008300781e-02,2.906040288507938385e-02,-1.018029823899269104e-01,5.357018858194351196e-02,4.841879382729530334e-02,-2.399152219295501709e-01,3.080863952636718750e-01,-2.472282052040100098e-01,-5.924335122108459473e-02,3.529893932864069939e-03,4.914423823356628418e-02,-1.018783226609230042e-01,-9.140267968177795410e-02,-6.821420043706893921e-02,3.727219626307487488e-02,-2.346913218498229980e-01,3.075305521488189697e-01,1.349108368158340454e-01,-1.341476142406463623e-01,1.573688834905624390e-01,3.602253273129463196e-02,3.827838599681854248e-01,-1.745749115943908691e-01,6.336758136749267578e-01,4.382032454013824463e-01,-4.363486915826797485e-02,1.654023528099060059e-01,-2.497493103146553040e-02,-2.442323230206966400e-02,-9.507476538419723511e-02,2.475168742239475250e-02,-3.665302395820617676e-01,-1.454804390668869019e-01,-3.225041627883911133e-01,8.177345991134643555e-02,2.314988970756530762e-01,4.994299113750457764e-01,1.633587479591369629e-01,2.621903121471405029e-01,-8.750110864639282227e-03,-1.623129844665527344e-01,3.249768316745758057e-01,1.792649775743484497e-01,-2.340880967676639557e-02,9.833842515945434570e-02,1.264463365077972412e-01,3.766472041606903076e-01,5.043060779571533203e-01,6.933655738830566406e-01,5.457080006599426270e-01,4.933836758136749268e-01,3.864742815494537354e-01,3.896686732769012451e-01,1.969470381736755371e-01,1.032048687338829041e-01,-1.403466314077377319e-01,-1.251981593668460846e-03,-9.028897434473037720e-02,8.740556240081787109e-02,-5.082302168011665344e-02,1.739999353885650635e-01,-9.087904542684555054e-02,1.540226936340332031e-01,-1.849243789911270142e-01,-1.166499964892864227e-02,2.228264696896076202e-03,1.974864155054092407e-01,-3.246231004595756531e-02,1.644202321767807007e-01,1.140366122126579285e-01,1.239080950617790222e-01,2.202164828777313232e-01,2.002957016229629517e-01,1.604662090539932251e-01,3.282775878906250000e-01,2.824743688106536865e-01,2.332290858030319214e-01,4.849811643362045288e-02,3.025672435760498047e-01,1.087647527456283569e-01,-2.374247834086418152e-02,4.578008875250816345e-02,-7.734116911888122559e-02,1.435022950172424316e-01,-2.037636041641235352e-01,-3.121909126639366150e-02,6.989226490259170532e-02,1.186490729451179504e-01,8.420057594776153564e-02,2.421660581603646278e-03,4.696421325206756592e-03,-3.255507349967956543e-02,3.311477228999137878e-02,-1.900814101099967957e-02,6.540261209011077881e-02,2.036921530961990356e-01,-8.160351961851119995e-02,1.240523979067802429e-01,1.047618091106414795e-01,2.174081057310104370e-01,1.900397390127182007e-01,-8.641169965267181396e-02,7.351988554000854492e-02,5.867522209882736206e-02,2.015284597873687744e-01,2.480605691671371460e-01,-9.663890302181243896e-02,3.069701194763183594e-01,8.548272401094436646e-02,2.094300091266632080e-01,1.323162764310836792e-01,1.173839643597602844e-01,1.993487328290939331e-01,-8.515716530382633209e-03,1.147290840744972229e-01,-2.213513851165771484e-02,1.015517935156822205e-01,1.308008879423141479e-01,2.427138835191726685e-01,1.468778401613235474e-01,8.631505072116851807e-03,2.022117562592029572e-02,7.532697916030883789e-02,5.393003299832344055e-02,1.457910537719726562e-01,-1.792823374271392822e-01,2.038727551698684692e-01,-4.309149517212063074e-04,7.625266443938016891e-03,2.521854937076568604e-01,1.272008419036865234e-01,1.952635347843170166e-01,-1.163743361830711365e-01,1.793492585420608521e-01,2.253997139632701874e-02,-1.396604776382446289e-01,1.668117344379425049e-01,-2.521508932113647461e-01,2.637263834476470947e-01,-1.075998768210411072e-01,1.634059846401214600e-01,4.209144040942192078e-02,2.201486378908157349e-01,2.106802016496658325e-01,1.872080117464065552e-01,8.742655068635940552e-02,1.339690089225769043e-01,1.316167414188385010e-01,2.793703079223632812e-01,6.318835914134979248e-02,1.581396460533142090e-01,3.472394347190856934e-01,1.752851903438568115e-01,5.145517364144325256e-02,1.626305282115936279e-01,-5.664709210395812988e-02,1.768629699945449829e-01,3.067570552229881287e-02,3.619053587317466736e-02,-9.443052858114242554e-02,-1.970933675765991211e-01,-1.299661695957183838e-01,-2.052543312311172485e-01,-4.539014771580696106e-02,-3.392856419086456299e-01,-2.505169808864593506e-01,-5.958970785140991211e-01,-5.433236956596374512e-01,-6.757769733667373657e-02,-6.167978793382644653e-02,-5.160158872604370117e-02,3.356191813945770264e-01,3.579602539539337158e-01,1.941171735525131226e-01,-6.195660680532455444e-02,5.225554481148719788e-02,1.763600856065750122e-01,-9.199210256338119507e-02,1.466574668884277344e-01,-3.006360307335853577e-02,-8.260319381952285767e-02,-4.550798609852790833e-02,-1.948628127574920654e-01,-2.151329815387725830e-02,-2.726104259490966797e-01,-2.598754465579986572e-01,-9.812887012958526611e-02,-2.002151906490325928e-01,-7.972714304924011230e-02,-8.171458542346954346e-02,-2.917539477348327637e-01,-3.343160450458526611e-01,-6.396834552288055420e-02,-1.205657273530960083e-01,-2.006701976060867310e-01,-9.704504162073135376e-02,-2.662470340728759766e-01,-1.795307993888854980e-01,-1.128808781504631042e-02,-2.760598063468933105e-01,-3.196404129266738892e-02,-1.954487562179565430e-01,-1.770293153822422028e-02,-9.468080103397369385e-02,-9.899703413248062134e-02,1.195527315139770508e-01,-1.070432439446449280e-01,-1.868489384651184082e-01,-7.982997223734855652e-03,4.704520106315612793e-02,-6.626465171575546265e-02,-1.201128065586090088e-01,-1.296261847019195557e-01,-1.180759742856025696e-01,-6.366629898548126221e-02,4.630334209650754929e-03,1.256527304649353027e-01,1.467499732971191406e-01,-3.439112333580851555e-04,-1.699746996164321899e-01,1.288965940475463867e-01,-6.699283141642808914e-03,9.283918887376785278e-02,-1.494404673576354980e-02,-1.011932268738746643e-03,1.449841558933258057e-01,1.613850444555282593e-01,2.010243684053421021e-01,1.367246955633163452e-01,1.532678306102752686e-01,-1.267800480127334595e-01,9.110566973686218262e-02,1.142581179738044739e-01,-1.700081378221511841e-01,-9.083208627998828888e-03,1.137482747435569763e-01,1.508615761995315552e-01,-5.408199131488800049e-02,1.283942312002182007e-01,7.545083761215209961e-02,-8.553203940391540527e-02,6.149076297879219055e-02,1.173660829663276672e-01,-2.344755828380584717e-01,1.634073406457901001e-01,6.188099831342697144e-02,1.066978052258491516e-01,4.006842151284217834e-02,-2.240373939275741577e-02,-4.215738549828529358e-02,2.825548052787780762e-01,1.466802805662155151e-01,1.105668917298316956e-01,-1.651368290185928345e-02,1.188554167747497559e-01,3.288356959819793701e-02,1.995637416839599609e-01,2.450135052204132080e-01,2.462515681982040405e-01,1.706076860427856445e-01,1.963631659746170044e-01,1.825316101312637329e-01,1.180866453796625137e-02,-1.733207143843173981e-02,1.738826930522918701e-01,-1.254608761519193649e-02,5.426232144236564636e-02,1.103315502405166626e-01,2.430720031261444092e-01,2.806808948516845703e-01,2.441507875919342041e-01,3.296599984169006348e-01,1.291851252317428589e-01,2.250366210937500000e-01,1.869978941977024078e-02,2.060850262641906738e-01,2.590595483779907227e-01,-2.138025127351284027e-02,2.545615732669830322e-01,-1.552529931068420410e-01,1.723461747169494629e-01,1.736114546656608582e-02,-2.112882584333419800e-01,2.459818124771118164e-01,-1.223125122487545013e-02,1.652079820632934570e-01,4.637175798416137695e-02,1.261118501424789429e-01,-3.418871760368347168e-01,-1.736644655466079712e-01,6.041649356484413147e-02,-8.025943487882614136e-02,-2.453791052103042603e-01,-5.245862603187561035e-01,-6.491080522537231445e-01,-6.287286281585693359e-01,-4.630112648010253906e-01,1.003754511475563049e-01,3.895644843578338623e-01,-4.985226988792419434e-01,3.113757967948913574e-01,-1.024849563837051392e-01,1.717985421419143677e-01,-1.745049059391021729e-01,3.631120175123214722e-02,3.308861553668975830e-01,2.976612746715545654e-01,5.844030380249023438e-01,4.015144109725952148e-01,3.552768826484680176e-01,3.296500146389007568e-01,1.258426606655120850e-01,9.376905858516693115e-02,6.770354509353637695e-02,3.469552695751190186e-01,3.328467905521392822e-02,9.348813444375991821e-02,1.237478181719779968e-01,-1.260541379451751709e-01,9.917128831148147583e-02,1.580283641815185547e-01,-6.117571517825126648e-02,1.405742764472961426e-01,-6.174173951148986816e-02,-9.327396005392074585e-02,1.678238213062286377e-01,-3.742452245205640793e-03,-2.455704212188720703e-01,-2.086653709411621094e-01,6.338869035243988037e-02,-2.375825196504592896e-01,7.335297018289566040e-02,-1.823571622371673584e-01,-2.429282516241073608e-01,-1.479599177837371826e-01,-7.776443660259246826e-02,-3.100043721497058868e-02,-3.605065047740936279e-01,7.104212790727615356e-02,-7.033132761716842651e-02,-1.303143799304962158e-01,-2.987981438636779785e-01,-1.796680539846420288e-01,-3.143789470195770264e-01,-1.593832224607467651e-01,-2.522590160369873047e-01,-3.385488390922546387e-01,-2.081451117992401123e-01,-2.001705616712570190e-01,-8.936768770217895508e-02,-2.436533421277999878e-01,-1.446970105171203613e-01,-2.033755481243133545e-01,-2.321061491966247559e-01,-2.382811754941940308e-01,-5.722391605377197266e-02,-6.889210548251867294e-03,-2.728121876716613770e-01,8.795142918825149536e-02,-9.426765888929367065e-02,-1.672883629798889160e-01,1.007510498166084290e-01,-1.734953671693801880e-01,-7.624514400959014893e-02,5.562783777713775635e-02,-2.261677086353302002e-01,-1.993048191070556641e-01,-1.277291923761367798e-01,-1.018084287643432617e-01,-2.996165752410888672e-01,6.644216366112232208e-03,1.476065516471862793e-01,-1.723688542842864990e-01,1.863213479518890381e-01,-2.215566299855709076e-02,-1.564820483326911926e-02,-7.656636834144592285e-02,1.110030934214591980e-01,2.018339335918426514e-01,2.164504826068878174e-01,-9.377297759056091309e-02,2.740258350968360901e-02,-3.879480808973312378e-02,3.326238095760345459e-01,5.907879397273063660e-02,1.057623028755187988e-01,2.747122645378112793e-01,1.350298523902893066e-02,1.934025883674621582e-01,1.365759819746017456e-01,-1.438447833061218262e-01,-9.436507523059844971e-02,1.657227128744125366e-01,9.077680855989456177e-02,-2.608461119234561920e-02,2.216590791940689087e-01,1.208485662937164307e-01,1.679932922124862671e-01,2.725499682128429413e-02,2.501056194305419922e-01,-9.268451482057571411e-02,2.743598222732543945e-01,5.491207912564277649e-02,2.877786755561828613e-01,-7.977854460477828979e-02,-9.873591363430023193e-02,-9.791193157434463501e-02,1.677486002445220947e-01,-3.826365619897842407e-02,7.005745172500610352e-02,-1.456663757562637329e-01,1.692977733910083771e-02,-8.936931192874908447e-02,-9.550484269857406616e-02,-3.700855746865272522e-02,-1.700428724288940430e-01,-9.553499519824981689e-02,-4.813472740352153778e-03,-5.006343498826026917e-02,1.205441728234291077e-01,-2.402378469705581665e-01,-1.087291836738586426e-01,-5.810059905052185059e-01,-1.197905912995338440e-01,-5.919715762138366699e-01,-3.445016443729400635e-01,5.063694715499877930e-01,2.324425280094146729e-01,3.163659572601318359e-01,-1.156620755791664124e-01,2.016805112361907959e-01,1.331125050783157349e-01,-2.366727963089942932e-02,-2.481587976217269897e-02,-1.456787586212158203e-01,-2.497764229774475098e-01,-1.390208005905151367e-01,-2.278267443180084229e-01,-1.529498770833015442e-02,-1.253886967897415161e-01,-8.342806994915008545e-02,-2.126801013946533203e-01,-9.878705441951751709e-02,7.614103704690933228e-02,-1.136554107069969177e-01,-4.151961952447891235e-02,-2.515554428100585938e-01,-5.233970880508422852e-01,-2.086290158331394196e-02,1.222681626677513123e-01,-1.744523271918296814e-02,-5.858611315488815308e-02,-2.539446055889129639e-01,-2.756597101688385010e-01,-7.728879153728485107e-02,5.642790719866752625e-02,5.981535091996192932e-02,-3.049438297748565674e-01,1.540569216012954712e-02,-3.384358063340187073e-02,1.574942283332347870e-02,5.891593545675277710e-02,9.379589557647705078e-02,2.738231606781482697e-02,1.472086906433105469e-01,-1.226881369948387146e-01,1.746443361043930054e-01,7.230751216411590576e-02,1.130222529172897339e-01,-2.346925437450408936e-01,1.821981370449066162e-01,-7.857216149568557739e-02,9.069850295782089233e-02,-3.939262777566909790e-02,8.267095685005187988e-02,-1.268357783555984497e-01,-1.406590491533279419e-01,9.967619925737380981e-02,-1.239471733570098877e-01,-1.057212874293327332e-01,-1.259565949440002441e-01,2.057791873812675476e-02,2.046482115983963013e-01,-3.434678614139556885e-01,-1.055263653397560120e-01,-2.174955010414123535e-01,-5.653803050518035889e-02,-1.718957573175430298e-01,-7.335387915372848511e-02,3.030677791684865952e-03,-2.428562194108963013e-01,-1.620812416076660156e-01,-1.252830326557159424e-01,-2.208880931138992310e-01,3.220244497060775757e-02,-2.436202317476272583e-01,-1.110069081187248230e-01,-2.924277186393737793e-01,-7.074303179979324341e-02,-1.928961426019668579e-01,1.710604429244995117e-01,-3.369787633419036865e-01,7.247257977724075317e-02,-1.794685721397399902e-01,-3.193362951278686523e-01,-3.451611995697021484e-01,-1.495336592197418213e-01,-7.006306946277618408e-02,-2.395810484886169434e-01,-3.965849578380584717e-01,-1.494739055633544922e-01,3.904401510953903198e-02,-3.361644148826599121e-01,-8.906516432762145996e-02,-1.177896112203598022e-01,-6.482195854187011719e-02,-2.107904702425003052e-01,1.189722493290901184e-01,-1.689103245735168457e-01,-5.477171018719673157e-02,-2.875213027000427246e-01,1.258808560669422150e-02,8.391575887799263000e-03,-6.290096044540405273e-02,5.495614558458328247e-02,6.569943577051162720e-02,1.244055666029453278e-02,3.256855309009552002e-01,-7.008019089698791504e-02,9.407955408096313477e-02,-4.149334039539098740e-03,-2.952374331653118134e-02,1.037191748619079590e-01,8.762104064226150513e-02,-3.489901125431060791e-01,1.042986884713172913e-01,1.078817620873451233e-01,7.911247014999389648e-02,-2.553505450487136841e-02,-1.038017049431800842e-01,-1.118268743157386780e-01,-7.629194110631942749e-02,-1.790132224559783936e-01,6.816270947456359863e-02,-3.877887725830078125e-01,-1.079048067331314087e-01,8.881016820669174194e-02,5.787578597664833069e-02,2.351800501346588135e-01,3.194087371230125427e-02,-1.365090310573577881e-01,-2.389923483133316040e-01,-1.431670337915420532e-01,1.625051051378250122e-01,2.470092028379440308e-01,-1.760680228471755981e-01,2.146905660629272461e-01,3.578656585887074471e-03,-2.624016404151916504e-01,4.811448156833648682e-01,7.080321311950683594e-01,2.399649769067764282e-01,4.846134781837463379e-01,1.883105635643005371e-01,-1.483039706945419312e-01,-4.583863019943237305e-01,-2.530335783958435059e-01,-3.084601163864135742e-01,2.244467474520206451e-02,7.487130910158157349e-02,6.541102379560470581e-02,1.707869172096252441e-01,-1.301468759775161743e-01,1.549488753080368042e-01,-1.327192634344100952e-01,1.273616552352905273e-01,-2.353077977895736694e-01,-1.406801640987396240e-01,-3.630204871296882629e-02,-1.493852138519287109e-01,-7.454747706651687622e-02,-8.369596302509307861e-02,7.083144783973693848e-02,-9.522286057472229004e-02,-2.179199270904064178e-02,-7.421673834323883057e-02,1.067924723029136658e-01,-3.431266844272613525e-01,4.103791713714599609e-01,-3.147362172603607178e-01,-1.962071210145950317e-01,5.407677590847015381e-02,1.052887812256813049e-01,-5.863365903496742249e-02,-1.956754922866821289e-01,-9.021139144897460938e-02,2.092821896076202393e-01,-4.082291573286056519e-02,2.204093486070632935e-01,-1.408871859312057495e-01,1.307462900876998901e-01,7.036843895912170410e-02,-1.186780408024787903e-01,-2.502006888389587402e-01,1.441930383443832397e-01,-2.075327485799789429e-01,1.877803057432174683e-01,-2.834182083606719971e-01,2.526341378688812256e-01,-1.577787101268768311e-01,-2.299987077713012695e-01,-6.505499035120010376e-02,4.541312903165817261e-02,1.042483821511268616e-01,-5.795083008706569672e-03,2.084084451198577881e-01,6.495510041713714600e-02,-2.109923213720321655e-02,-2.837538719177246094e-02,2.381629943847656250e-01,3.257825970649719238e-01,-2.000425755977630615e-02,-2.240263372659683228e-01,1.735004931688308716e-01,-9.036562591791152954e-02,-1.978688538074493408e-01,-9.871514886617660522e-02,-1.394356042146682739e-01,-2.466534972190856934e-01,-1.029685884714126587e-02,-2.594599127769470215e-01,3.170399069786071777e-01,-2.123339623212814331e-01,3.620237857103347778e-02,-2.164308279752731323e-01,-1.811876296997070312e-01,-3.468489646911621094e-02,-2.412587702274322510e-01,8.537673950195312500e-02,4.949006065726280212e-02,-1.386406421661376953e-01,-3.494636621326208115e-03,-9.241825342178344727e-02,1.392061263322830200e-01,-1.802473664283752441e-01,1.006438136100769043e-01,-1.307236868888139725e-02,-9.725234471261501312e-03,2.887504547834396362e-02,-5.418427661061286926e-02,-1.288681942969560623e-02,-1.411723997443914413e-02,4.337868690490722656e-01,5.584229715168476105e-03,1.574174910783767700e-01,-2.105747722089290619e-02,1.096426844596862793e-01,1.179036572575569153e-01,4.226117581129074097e-02,-2.279190272092819214e-01,7.000082731246948242e-02,-3.593365475535392761e-02,-8.499206602573394775e-02,-2.297105193138122559e-01,2.601494193077087402e-01,5.186723545193672180e-03,1.446166336536407471e-01,-1.347863487899303436e-02,1.017178408801555634e-02,-4.561930149793624878e-02,1.832197606563568115e-01,-9.491922706365585327e-02,-1.344285011291503906e-01,-2.849436104297637939e-01,-1.829155385494232178e-01,-1.065856963396072388e-01,6.130409836769104004e-01,9.329702854156494141e-01,3.115156292915344238e-01,7.675459235906600952e-02,-1.321080625057220459e-01,4.137800633907318115e-01,1.439001969993114471e-02,4.822256416082382202e-02,1.857690662145614624e-01,1.025150567293167114e-01,-2.065267264842987061e-01,3.872666060924530029e-01,2.097078561782836914e-01,-7.095654010772705078e-01,-5.623558908700942993e-02,5.270804464817047119e-02,-7.180209457874298096e-02,-7.288300991058349609e-02,5.812708660960197449e-02,-1.239221990108489990e-01,-2.103203162550926208e-02,1.382329314947128296e-01,-6.552041321992874146e-02,8.889376372098922729e-02,-1.053438894450664520e-02,1.163801550865173340e-01,6.991709768772125244e-02,1.332594305276870728e-01,6.940253823995590210e-02,-2.521897666156291962e-02,9.809273481369018555e-02,1.769231110811233521e-01,-1.060476973652839661e-01,1.140064522624015808e-01,-1.769754453562200069e-04,9.102053195238113403e-02,9.795866906642913818e-02,2.543973550200462341e-02,7.527913898229598999e-02,-6.200641393661499023e-02,-7.880918681621551514e-03,4.430886730551719666e-02,1.700561307370662689e-02,9.236203134059906006e-02,-1.055234223604202271e-01,1.108458545058965683e-02,-1.611445099115371704e-01,5.541330948472023010e-02,-1.276768147945404053e-01,-7.172488421201705933e-02,6.176578626036643982e-02,-1.544391363859176636e-01,-9.128613770008087158e-02,-1.809755340218544006e-02,4.588616266846656799e-02,-1.002273783087730408e-01,6.441457569599151611e-02,-5.428345873951911926e-02,-7.514010369777679443e-02,4.014725238084793091e-02,-9.172589518129825592e-03,-4.764613136649131775e-02,7.035229820758104324e-03,-1.363576054573059082e-01,1.831305772066116333e-01,-2.186478488147258759e-02,-1.390643138438463211e-02,3.973678499460220337e-02,-1.077298074960708618e-01,7.636333256959915161e-02,2.536891959607601166e-02,6.223319470882415771e-02,5.242991726845502853e-03,1.129612103104591370e-01,5.069209262728691101e-02,1.417695730924606323e-01,-7.013024296611547470e-03,2.007835954427719116e-01,-5.362061411142349243e-02,1.154154688119888306e-01,2.240343093872070312e-01,-2.972787246108055115e-02,-1.102412212640047073e-02,1.712045446038246155e-02,7.058691978454589844e-02,1.832910478115081787e-01,3.204152733087539673e-02,-5.701253656297922134e-03,1.497419327497482300e-01,1.180167943239212036e-01,-9.886542707681655884e-02,1.375758498907089233e-01,1.022401377558708191e-01,-8.977207541465759277e-02,1.881467700004577637e-01,2.655670233070850372e-02,-7.109199650585651398e-04,1.167460307478904724e-01,4.433673992753028870e-02,8.023178088478744030e-04,1.340596377849578857e-01,-1.109893396496772766e-01,1.496334075927734375e-01,8.561257272958755493e-02,6.917206197977066040e-02,1.825391873717308044e-02,1.354765743017196655e-01,2.580748312175273895e-02,5.189325287938117981e-02,7.358117401599884033e-02,8.386746048927307129e-03,2.124476730823516846e-01,9.927543252706527710e-02,9.947534650564193726e-02,4.996046051383018494e-02,1.064117029309272766e-01,-6.087327748537063599e-02,1.559334248304367065e-01,1.247244179248809814e-01,1.420401632785797119e-01,-1.443285644054412842e-01,2.623742520809173584e-01,1.777875721454620361e-01,-1.056488305330276489e-01,2.683912217617034912e-01,1.991516798734664917e-01,-1.003391295671463013e-01,-5.021475628018379211e-02,-1.496510356664657593e-01,-8.087346553802490234e-01,8.941592574119567871e-01,9.730316996574401855e-01,-5.733057856559753418e-01,2.305645495653152466e-01,-9.634578973054885864e-02,-1.364528834819793701e-01,-1.431219726800918579e-01,4.119434654712677002e-01,8.790075778961181641e-01,5.062907934188842773e-01,2.025506645441055298e-01,-3.949516713619232178e-01,-8.421409875154495239e-02,-1.104586496949195862e-01,-6.602083146572113037e-02,-3.299083113670349121e-01,-6.018662452697753906e-02,-1.254248023033142090e-01,-9.518993645906448364e-02,6.189121678471565247e-02,2.738413400948047638e-02,-1.740454286336898804e-01,1.417679190635681152e-01,1.257839798927307129e-01,-2.517140805721282959e-01,3.862609341740608215e-02,6.403315812349319458e-02,6.134873628616333008e-02,-6.129298731684684753e-02,6.882454454898834229e-02,-4.522890225052833557e-02,2.081110477447509766e-01,2.136070728302001953e-01,-8.130349963903427124e-02,8.394598215818405151e-02,-8.656080812215805054e-02,1.609418541193008423e-01,-2.320489287376403809e-02,1.135844662785530090e-01,1.026860717684030533e-02,8.344439417123794556e-02,-1.123305261135101318e-01,1.504881959408521652e-02,-1.096317544579505920e-01,4.178014397621154785e-02,2.923843264579772949e-02,1.437850482761859894e-02,-5.239613354206085205e-02,-1.506582945585250854e-01,-1.300022304058074951e-01,-2.096042633056640625e-01,4.376219213008880615e-01,-1.535412818193435669e-01,-4.962317645549774170e-02,1.492830812931060791e-01,-7.889264076948165894e-02,-6.938111782073974609e-02,-3.756646215915679932e-01,-6.599643081426620483e-02,7.635895628482103348e-03,-1.621390581130981445e-01,-2.703000605106353760e-01,8.505775034427642822e-02,-8.441202342510223389e-03,-1.423638127744197845e-02,-1.456564962863922119e-01,-2.412903159856796265e-01,2.011392638087272644e-02,-2.439992874860763550e-01,-1.238789185881614685e-01,-1.824040859937667847e-01,-1.217488348484039307e-01,-3.233631849288940430e-01,-1.332037895917892456e-01,-1.202691495418548584e-01,-1.428522169589996338e-01,-1.411365419626235962e-01,-7.255284488201141357e-02,1.673868596553802490e-01,-8.340657502412796021e-02,-2.008694559335708618e-01,-3.916796743869781494e-01,8.882983028888702393e-02,-2.500766515731811523e-01,1.628447473049163818e-01,-3.143786489963531494e-01,-2.140186727046966553e-03,1.441617310047149658e-01,-4.859381020069122314e-01,8.846591413021087646e-02,-1.724144220352172852e-01,-5.218828096985816956e-02,-7.788731902837753296e-02,2.972124703228473663e-02,-3.719406202435493469e-02,5.138718709349632263e-02,-5.200755968689918518e-02,-1.125891134142875671e-01,8.890494704246520996e-02,1.445953175425529480e-02,-1.220047175884246826e-01,4.926698654890060425e-02,9.592414647340774536e-02,2.273587733507156372e-01,2.473151087760925293e-01,1.369054466485977173e-01,9.260289371013641357e-03,3.287266194820404053e-02,-3.283459320664405823e-02,2.796480953693389893e-01,1.485611945390701294e-01,1.826096475124359131e-01,1.927845925092697144e-01,-4.224105924367904663e-02,9.432930499315261841e-02,5.538607761263847351e-02,-9.071175754070281982e-02,1.192776188254356384e-01,1.404828876256942749e-01,2.371050566434860229e-01,2.348300516605377197e-01,-1.205567177385091782e-02,3.681471943855285645e-01,5.851840972900390625e-02,8.618059009313583374e-02,-4.618932008743286133e-01,-5.440952777862548828e-01,-7.192767262458801270e-01,-3.125435709953308105e-01,-5.509441345930099487e-02,6.499591469764709473e-01,3.196046948432922363e-01,-8.983852714300155640e-02,3.436372876167297363e-01,2.710044085979461670e-01,4.332549571990966797e-01,3.374551236629486084e-01,5.283138155937194824e-01,2.761394679546356201e-01,1.775339990854263306e-01,2.872644960880279541e-01,-1.977011710405349731e-01,-3.049671351909637451e-01,4.331878572702407837e-02,6.551808118820190430e-02,1.064983978867530823e-01,-4.160121083259582520e-02,7.722064107656478882e-02,-3.208813723176717758e-04,-1.095949634909629822e-01,5.960444733500480652e-02,-5.053345859050750732e-02,-1.673342734575271606e-01,1.965887397527694702e-01,3.903421387076377869e-02,1.778116971254348755e-01,-6.957384198904037476e-02,-5.713837221264839172e-02,-1.597742438316345215e-01,2.281539589166641235e-01,-1.955228149890899658e-01,1.878642141819000244e-01,-1.424240767955780029e-01,-1.069805249571800232e-01,1.413525640964508057e-01,-3.256631270051002502e-02,-6.252710521221160889e-02,4.367210343480110168e-02,5.003963038325309753e-02,8.213360607624053955e-02,1.645730137825012207e-01,1.393994688987731934e-01,2.047347463667392731e-02,2.554084733128547668e-02,3.253200948238372803e-01,1.141900122165679932e-01,-2.281163074076175690e-02,1.573081165552139282e-01,-5.232746526598930359e-02,4.165734946727752686e-01,6.823610514402389526e-02,5.137951672077178955e-02,6.862518936395645142e-02,2.295273542404174805e-01,-6.453210115432739258e-02,-4.353107139468193054e-02,1.153966411948204041e-01,-8.054634183645248413e-02,1.844141334295272827e-01,-1.325100660324096680e-01,2.390328943729400635e-01,7.922621443867683411e-04,9.825323522090911865e-02,1.538009494543075562e-01,-2.290170267224311829e-02,2.647481299936771393e-02,4.055266454815864563e-02,3.297341167926788330e-01,2.089283079840242863e-04,1.606621444225311279e-01,5.985342711210250854e-02,1.053254082798957825e-01,2.882541157305240631e-02,-3.270325437188148499e-02,3.090335428714752197e-01,3.093130327761173248e-02,2.597033679485321045e-01,9.686600416898727417e-02,2.038657963275909424e-01,2.521918714046478271e-01,-7.421418279409408569e-02,2.098122984170913696e-01,9.158050268888473511e-02,-2.363770455121994019e-02,1.968098878860473633e-01,1.675111949443817139e-01,6.581951677799224854e-02,2.941457927227020264e-01,9.815978258848190308e-02,3.564550280570983887e-01,2.481961250305175781e-01,-1.337261684238910675e-02,4.960916340351104736e-01,3.173148036003112793e-01,3.310451209545135498e-01,2.203420251607894897e-01,3.846202790737152100e-01,3.058434724807739258e-01,4.005178809165954590e-01,2.773869931697845459e-01,2.072009593248367310e-01,1.950713247060775757e-01,3.324449360370635986e-01,3.683801293373107910e-01,8.271329104900360107e-02,2.368212789297103882e-01,1.375193148851394653e-01,2.388634681701660156e-01,6.691581010818481445e-02,3.052278757095336914e-01,-1.166958659887313843e-01,-1.123888138681650162e-02,1.812116056680679321e-02,1.894533336162567139e-01,1.665661782026290894e-01,-8.872158080339431763e-02,-1.332205384969711304e-01,-1.140454690903425217e-02,-8.366177976131439209e-02,-1.541272401809692383e-01,-1.647073030471801758e-01,-5.052783340215682983e-02,1.015827711671590805e-02,-5.737154185771942139e-02,8.828946202993392944e-02,-4.931235611438751221e-01,-9.722413867712020874e-02,8.560806512832641602e-01,7.127120494842529297e-01,6.915953159332275391e-01,5.941748991608619690e-02,1.576541215181350708e-01,4.341672658920288086e-01,-1.465982198715209961e-01,1.321267485618591309e-01,5.324963331222534180e-01,8.815172910690307617e-01,6.853733062744140625e-01,2.125279605388641357e-01,3.778518363833427429e-02,-2.352431267499923706e-01,2.595306746661663055e-02,1.689338833093643188e-01,1.689549535512924194e-01,2.008293867111206055e-01,-5.288522318005561829e-02,2.456984072923660278e-01,1.253899484872817993e-01,1.486032903194427490e-01,2.276235073804855347e-02,-2.220418304204940796e-02,-5.576141923666000366e-02,-2.084148973226547241e-01,8.834058791399002075e-02,5.063233524560928345e-02,7.033689320087432861e-02,2.025560103356838226e-02,1.434984058141708374e-02,-4.717307537794113159e-02,1.916134655475616455e-01,-7.050815224647521973e-02,-1.310789734125137329e-01,-2.563527822494506836e-01,-2.166163623332977295e-01,1.371079981327056885e-01,-3.103668987751007080e-01,4.827875643968582153e-02,-2.101603299379348755e-01,-8.762308210134506226e-02,-1.213277578353881836e-01,2.288746833801269531e-02,1.413043588399887085e-01,1.002134829759597778e-01,-1.355137974023818970e-01,-5.156251415610313416e-02,-1.469481885433197021e-01,1.645727157592773438e-01,-2.104993462562561035e-01,1.523609161376953125e-01,1.609908491373062134e-01,-3.384814411401748657e-02,5.925309285521507263e-02,-1.643115133047103882e-01,4.658169299364089966e-02,-3.801333010196685791e-01,1.587828993797302246e-01,1.510416716337203979e-01,1.238184347748756409e-01,3.259984403848648071e-02,-1.820932924747467041e-01,1.105284020304679871e-01,-1.803802400827407837e-01,2.009883224964141846e-01,1.188911274075508118e-01,6.050353497266769409e-02,-4.012382030487060547e-02,-2.032784745097160339e-02,-1.641113013029098511e-01,2.383109480142593384e-01,-8.283155038952827454e-03,8.712051808834075928e-02,-9.766662120819091797e-02,-2.236680239439010620e-01,1.809047013521194458e-01,-1.738304458558559418e-02,3.304090723395347595e-02,2.452575415372848511e-01,-1.058140024542808533e-01,-1.115250438451766968e-01,1.768601983785629272e-01,8.694858849048614502e-02,2.428832277655601501e-02,3.453896939754486084e-02,1.457745730876922607e-01,-1.223241835832595825e-01,-1.154460608959197998e-01,-1.058522611856460571e-01,-4.224172607064247131e-02,-1.339587718248367310e-01,-9.818932414054870605e-02,-1.558194607496261597e-01,-1.925832405686378479e-02,-1.814788579940795898e-01,-1.256802976131439209e-01,9.922410547733306885e-02,-2.270406037569046021e-01,-1.528113335371017456e-01,9.541878849267959595e-02,-3.111851401627063751e-02,-1.076476424932479858e-01,7.232300937175750732e-02,5.214909836649894714e-02,1.731977909803390503e-01,-2.955510467290878296e-02,-2.541939355432987213e-02,7.212822139263153076e-02,2.553703486919403076e-01,7.918720692396163940e-02,1.195363104343414307e-01,-1.461185812950134277e-01,-4.436982423067092896e-02,2.377418279647827148e-01,3.017556481063365936e-02,3.583045005798339844e-01,4.790866002440452576e-02,2.002516686916351318e-01,5.356572219170629978e-04,4.204995334148406982e-01,3.628668189048767090e-01,4.831485450267791748e-01,3.062861263751983643e-01,8.383332751691341400e-03,5.097850412130355835e-02,1.606671363115310669e-01,1.461646705865859985e-01,4.348569512367248535e-01,2.684293985366821289e-01,3.719363510608673096e-01,3.043795824050903320e-01,1.206565797328948975e-01,1.870981305837631226e-01,3.526135161519050598e-02,3.305254876613616943e-01,-5.832447484135627747e-02,-7.824591398239135742e-01,-2.700983881950378418e-01,2.086145132780075073e-01,-1.964563727378845215e-01,-1.609586626291275024e-01,1.273320317268371582e-01,1.368562579154968262e-01,1.037563085556030273e-01,2.040986269712448120e-01,1.874696165323257446e-01,-8.659363724291324615e-03,2.391356080770492554e-01,-6.129911541938781738e-02,-6.498850882053375244e-02,3.876778483390808105e-02,6.798293441534042358e-02,2.979879826307296753e-02,-4.728570953011512756e-02,3.950972482562065125e-02,-5.376313254237174988e-02,-1.026053130626678467e-01,8.333107456564903259e-03,-6.286483258008956909e-02,-1.081830710172653198e-01,-1.498214304447174072e-01,-4.743606224656105042e-02,-9.680339694023132324e-02,-1.008636057376861572e-01,6.568559259176254272e-02,-2.051898688077926636e-01,-2.363440208137035370e-02,-6.574481725692749023e-02,-1.556477546691894531e-01,1.452040970325469971e-01,-4.712904617190361023e-02,2.649086117744445801e-01,-7.221493870019912720e-02,2.098797410726547241e-01,-1.304329782724380493e-01,-7.478312402963638306e-02,4.921361687593162060e-04,-4.786653816699981689e-02,9.161023795604705811e-02,-8.536742627620697021e-02,4.449009522795677185e-02,3.598704934120178223e-01,1.224725879728794098e-02,5.597824696451425552e-03,8.061369508504867554e-02,-6.061942502856254578e-02,3.336396440863609314e-02,-1.299059540033340454e-01,1.551530808210372925e-01,-2.596979439258575439e-01,2.065037786960601807e-01,-1.964722275733947754e-01,2.170441299676895142e-02,1.188419908285140991e-01,-2.503253519535064697e-01,1.311321258544921875e-01,9.907091967761516571e-03,-1.747992187738418579e-01,3.760958462953567505e-02,-1.101929545402526855e-01,-1.262354105710983276e-01,2.027897834777832031e-01,-4.881078004837036133e-02,1.450522989034652710e-01,-1.440997272729873657e-01,8.210582286119461060e-02,-1.070824712514877319e-01,-1.071606501936912537e-01,7.042599469423294067e-02,2.053706645965576172e-01,1.085994765162467957e-01,-2.015892416238784790e-01,3.187616169452667236e-01,1.087532937526702881e-01,-2.796787023544311523e-02,1.869899034500122070e-02,1.443792581558227539e-01,1.645591706037521362e-01,-1.344895362854003906e-01,2.131914496421813965e-01,1.011824682354927063e-01,1.232120543718338013e-01,3.290195167064666748e-01,1.424851566553115845e-01,2.862720191478729248e-01,2.867767810821533203e-01,7.737869024276733398e-02,-2.069666981697082520e-02,2.442669309675693512e-02,2.094888091087341309e-01,7.953921705484390259e-02,-6.024207919836044312e-02,2.561956457793712616e-02,-5.797994881868362427e-02,2.683610841631889343e-02,-8.785189688205718994e-02,-2.653968147933483124e-02,1.470196439186111093e-04,-5.544972792267799377e-02,-1.725327372550964355e-01,7.849874347448348999e-02,-1.339586675167083740e-01,-2.375845313072204590e-01,4.773251339793205261e-02,-2.565058171749114990e-01,-2.339319698512554169e-02,-3.857088088989257812e-02,-2.198249101638793945e-02,-4.571138694882392883e-02,2.749943137168884277e-01,-3.654330223798751831e-02,-1.115910932421684265e-01,7.026475071907043457e-01,-1.375585049390792847e-01,-1.221168160438537598e+00,1.894573122262954712e-01,7.890816330909729004e-01,1.438485383987426758e-01,-5.515427514910697937e-02,1.088732779026031494e-01,2.974345386028289795e-01,1.777116805315017700e-01,2.373938411474227905e-01,5.449473857879638672e-01,1.764710396528244019e-01,2.234789915382862091e-02,-4.996138811111450195e-01,-6.392218470573425293e-01,-5.883192420005798340e-01,-3.137097954750061035e-01,2.278725951910018921e-01,2.349717728793621063e-02,2.297435104846954346e-01,-1.768178194761276245e-01,1.754893958568572998e-01,7.932269945740699768e-04,1.263783127069473267e-01,1.498250514268875122e-01,-1.389830708503723145e-01,-1.058172509074211121e-01,5.819690972566604614e-02,8.745791390538215637e-03,1.939349919557571411e-01,-6.088140886276960373e-03,-8.168490976095199585e-02,1.145912632346153259e-01,-1.201920956373214722e-01,1.575706750154495239e-01,-4.287057369947433472e-02,-2.997208535671234131e-01,-1.704442352056503296e-01,-2.345281392335891724e-01,-1.280997991561889648e-01,-1.995991021394729614e-01,-2.425460815429687500e-01,-2.887343764305114746e-01,-2.563250660896301270e-01,7.865797728300094604e-02,-1.651567071676254272e-01,-2.248289622366428375e-02,-1.357529163360595703e-01,-1.003316119313240051e-01,-1.209387648850679398e-02,-6.920385360717773438e-02,8.037766069173812866e-02,-1.435885876417160034e-01,2.074865102767944336e-01,-6.489923596382141113e-02,-1.166689246892929077e-01,-1.426972895860671997e-01,-1.481123417615890503e-01,1.663844436407089233e-01,-3.158922791481018066e-01,3.458913043141365051e-02,-1.060999482870101929e-01,9.376917034387588501e-02,-2.679903209209442139e-01,1.925719678401947021e-01,-1.057312265038490295e-01,-2.511497735977172852e-01,-4.356810823082923889e-02,-2.321300804615020752e-01,5.804159864783287048e-02,-2.377257794141769409e-01,9.068655967712402344e-02,-2.210885733366012573e-01,-9.080526232719421387e-02,-1.300181299448013306e-01,-7.345902174711227417e-02,-6.856810301542282104e-02,4.611745476722717285e-02,-1.178212761878967285e-01,7.148833572864532471e-02,1.280196607112884521e-01,-2.999260127544403076e-01,1.573995351791381836e-01,-1.262824684381484985e-01,-1.976283341646194458e-01,8.644569665193557739e-02,5.043224245309829712e-02,-8.519399166107177734e-02,-6.063947081565856934e-02,-4.625185579061508179e-02,-2.972031012177467346e-02,-1.098724007606506348e-01,1.485955268144607544e-01,4.342669621109962463e-02,2.030209265649318695e-02,-2.150742337107658386e-02,1.590426564216613770e-01,1.034585908055305481e-01,2.866469323635101318e-01,1.675756722688674927e-01,1.316117644309997559e-01,1.784381717443466187e-01,1.561020594090223312e-02,-2.692232131958007812e-01,1.236500963568687439e-02,2.269335323944687843e-03,-2.284945100545883179e-01,-4.581444896757602692e-03,1.596448272466659546e-01,-1.129466965794563293e-01,1.422595530748367310e-01,-1.483006477355957031e-01,-8.927652239799499512e-02,-6.999797374010086060e-02,-4.500205218791961670e-01,1.237614899873733521e-01,-5.461423471570014954e-02,-3.301302716135978699e-02,-4.056207835674285889e-02,2.081531099975109100e-02,1.257594823837280273e-01,1.550351828336715698e-01,3.334154486656188965e-01,3.278899565339088440e-02,4.205772653222084045e-02,2.904203534126281738e-01,9.013770818710327148e-01,1.031718492507934570e+00,9.888320565223693848e-01,2.668549120426177979e-01,-2.945642173290252686e-01,-4.339495897293090820e-01,1.613393053412437439e-02,3.600395321846008301e-01,-4.015098139643669128e-02,-2.067538946866989136e-01,-1.026062294840812683e-01,1.142880395054817200e-01,-4.270986840128898621e-02,1.084509044885635376e-01,5.018573999404907227e-01,5.484910011291503906e-01,3.555656075477600098e-01,-3.864061785861849785e-03,-6.447874009609222412e-02,-7.731638848781585693e-02,1.343405991792678833e-01,-1.013193726539611816e-01,-1.125135719776153564e-01,1.275551021099090576e-01,1.126940473914146423e-01,-2.291678264737129211e-02,4.392341896891593933e-02,-1.408296823501586914e-01,-4.329850897192955017e-02,-1.939885318279266357e-01,-1.227252483367919922e-01,-8.730733394622802734e-02,-1.159826442599296570e-01,-1.664412170648574829e-01,-2.281990349292755127e-01,-2.894289493560791016e-01,-1.110311225056648254e-01,-3.298444300889968872e-02,-2.312965691089630127e-01,1.689404547214508057e-01,-1.767095327377319336e-01,-1.497578620910644531e-01,1.509649679064750671e-02,8.905836381018161774e-03,2.525164484977722168e-01,1.490354686975479126e-01,7.981200516223907471e-02,3.251531720161437988e-02,-1.092480793595314026e-01,7.785466313362121582e-02,2.676698565483093262e-01,3.547411784529685974e-02,7.351701706647872925e-02,6.305529177188873291e-02,-2.008395344018936157e-01,-3.430874645709991455e-02,-1.523804515600204468e-01,4.188288748264312744e-02,5.846245959401130676e-02,-1.684250086545944214e-01,4.240555223077535629e-03,1.029202044010162354e-01,-1.924609094858169556e-01,-1.146627590060234070e-01,6.861516088247299194e-02,-6.535844504833221436e-02,1.144721359014511108e-01,5.488194292411208153e-04,1.721842139959335327e-01,-1.166385784745216370e-02,2.291037291288375854e-01,4.708993248641490936e-03,-4.584784433245658875e-02,-1.277195662260055542e-01,6.774102151393890381e-02,1.083597838878631592e-01,6.242031231522560120e-02,-6.625563651323318481e-02,2.176144160330295563e-03,1.823794469237327576e-02,-1.228822991251945496e-01,1.169747207313776016e-02,-7.853285060264170170e-04,7.673541456460952759e-02,5.090859532356262207e-02,2.697233855724334717e-01,-1.554813235998153687e-01,-8.188077062368392944e-02,-2.375834882259368896e-01,9.356094896793365479e-02,1.067677363753318787e-01,3.550127148628234863e-02,1.239641606807708740e-01,-6.153744831681251526e-02,-3.621540591120719910e-02,-2.051613628864288330e-01,-1.237906217575073242e-01,-1.530523896217346191e-01,9.131778031587600708e-02,-6.109441071748733521e-02,7.730773091316223145e-02,-1.854923740029335022e-02,-1.249471772462129593e-02,-1.505267620086669922e-01,-8.931659162044525146e-02,1.165273785591125488e-02,1.902223564684391022e-02,3.169834315776824951e-01,-3.856955096125602722e-02,8.136619627475738525e-02,-1.729132607579231262e-02,-1.075691655278205872e-01,1.049431860446929932e-01,2.496575862169265747e-01,6.212120503187179565e-02,8.754748851060867310e-02,6.624760478734970093e-02,2.934222519397735596e-01,1.642611324787139893e-01,1.494312286376953125e-01,2.243463695049285889e-01,-5.832813680171966553e-02,1.137575358152389526e-01,3.228794336318969727e-01,2.844419181346893311e-01,3.148006796836853027e-01,3.480480909347534180e-01,3.122805058956146240e-01,3.090232312679290771e-01,4.909169375896453857e-01,7.904134690761566162e-02,-6.702168583869934082e-01,-1.108555555343627930e+00,-8.141299486160278320e-01,-4.806591197848320007e-02,-1.013045106083154678e-02,4.042034745216369629e-01,3.480512201786041260e-01,5.768438577651977539e-01,4.344482123851776123e-01,4.668072462081909180e-01,6.321135163307189941e-02,-3.425320386886596680e-01,-3.950876593589782715e-01,-3.182865977287292480e-01,-2.029433697462081909e-01,-2.375715821981430054e-01,-1.135136187076568604e-02,-1.157536171376705170e-02,-4.050072282552719116e-02,4.922859743237495422e-02,-2.804146520793437958e-02,3.116231039166450500e-02,-1.748141795396804810e-01,3.852245956659317017e-02,-4.237023741006851196e-02,-1.371380127966403961e-02,-6.189325824379920959e-03,-9.080230444669723511e-02,1.897751986980438232e-01,-4.492670763283967972e-03,1.704604327678680420e-01,2.114327251911163330e-02,-9.530688822269439697e-02,-7.954563945531845093e-02,2.819380760192871094e-01,2.304616756737232208e-02,-1.741709560155868530e-02,1.421642452478408813e-01,4.004423320293426514e-02,-1.607097312808036804e-02,2.932053525000810623e-03,-7.189655676484107971e-03,-4.615275189280509949e-02,9.054782800376415253e-03,-1.878397166728973389e-02,1.096716895699501038e-01,-7.220797706395387650e-03,3.831444308161735535e-02,1.099610254168510437e-01,3.343426063656806946e-02,8.415349572896957397e-02,1.270959526300430298e-01,2.140577882528305054e-01,1.244142577052116394e-01,1.307559311389923096e-01,8.610411733388900757e-02,2.283596992492675781e-01,1.344917714595794678e-02,6.319702416658401489e-02,2.237340658903121948e-01,1.326212193816900253e-02,5.817949399352073669e-02,-2.657168544828891754e-03,2.384989559650421143e-01,1.731007695198059082e-01,-4.953277483582496643e-02,6.347163766622543335e-02,2.754948509391397238e-04,-4.189663752913475037e-02,1.246322467923164368e-01,1.158926337957382202e-01,1.649443060159683228e-01,1.409330666065216064e-01,1.880129054188728333e-02,1.553054451942443848e-01,1.356427073478698730e-01,-1.765827983617782593e-01,2.068301141262054443e-01,1.325932294130325317e-01,2.081698924303054810e-01,4.973633587360382080e-02,-1.303463429212570190e-01,3.029710054397583008e-01,-7.857075333595275879e-02,1.828808635473251343e-01,-4.649028927087783813e-02,9.204186499118804932e-02,1.499908138066530228e-02,-6.464911624789237976e-03,5.563377402722835541e-03,2.280625700950622559e-01,-1.423576381057500839e-02,1.110115423798561096e-01,8.729841560125350952e-02,3.765928000211715698e-02,4.535909369587898254e-02,-5.621669813990592957e-02,4.668256267905235291e-02,1.098032817244529724e-01,7.128529995679855347e-02,6.633970141410827637e-02,8.858443051576614380e-02,1.789949983358383179e-01,1.674408912658691406e-01,3.543178439140319824e-01,3.026338480412960052e-02,1.646231859922409058e-01,3.682601451873779297e-01,1.160530745983123779e-01,7.104621082544326782e-02,3.158685564994812012e-01,8.606496453285217285e-02,2.238572090864181519e-01,1.282401829957962036e-01,1.058601066470146179e-01,1.377752721309661865e-01,9.763058274984359741e-02,2.583962678909301758e-01,-4.958362132310867310e-02,4.283071495592594147e-03,2.614731788635253906e-01,3.042927756905555725e-02,6.868877972010523081e-05,4.430044069886207581e-02,2.473111003637313843e-01,6.019129231572151184e-02,7.220342755317687988e-02,-3.535904586315155029e-01,-6.729233860969543457e-01,-1.117731928825378418e+00,-4.442556798458099365e-01,6.501079201698303223e-01,3.784613609313964844e-01,7.954955101013183594e-02,2.806530594825744629e-01,-2.474922388792037964e-01,-1.205032318830490112e-01,4.567944109439849854e-01,8.192803263664245605e-01,7.296804189682006836e-01,4.708427786827087402e-01,3.399672508239746094e-01,6.639838963747024536e-02,2.643824554979801178e-02,-4.171658456325531006e-01,-4.947857186198234558e-02,-4.821717441082000732e-01,1.982978545129299164e-02,-1.026918962597846985e-01,8.853456377983093262e-02,-1.961721479892730713e-02,1.211398467421531677e-01,7.097149640321731567e-02,1.041220277547836304e-01,1.538964956998825073e-01,-6.618098914623260498e-02,-9.131281077861785889e-02,2.070603221654891968e-01,3.699623048305511475e-02,-9.467397816479206085e-03,7.401965558528900146e-02,-1.122165843844413757e-01,1.745113581418991089e-01,8.884857408702373505e-03,2.776147127151489258e-01,5.195128172636032104e-02,2.573811709880828857e-01,-2.780803143978118896e-01,1.208753064274787903e-01,1.632956117391586304e-01,-6.252560764551162720e-02,-7.556856423616409302e-02,-2.854334712028503418e-01,-1.398380547761917114e-01,-3.466034233570098877e-01,3.561627492308616638e-02,-5.068634822964668274e-02,1.226168870925903320e-01,-5.704364553093910217e-02,-1.130566373467445374e-01,6.021233275532722473e-02,-1.712654531002044678e-01,-2.365847229957580566e-01,-9.531904011964797974e-02,-2.889890782535076141e-02,-1.316202729940414429e-01,9.858432412147521973e-02,2.318086475133895874e-02,2.712159045040607452e-02,-1.878084391355514526e-01,4.483062773942947388e-03,-1.208871304988861084e-01,-2.778013646602630615e-01,-4.762845635414123535e-01,5.880923941731452942e-02,-3.746814280748367310e-02,-2.182139307260513306e-01,-1.840345934033393860e-02,-4.153514280915260315e-02,2.860044687986373901e-02,-3.462916985154151917e-02,-7.141354680061340332e-02,8.260954928118735552e-05,1.576014757156372070e-01,3.342083469033241272e-02,-3.723773360252380371e-01,1.410066634416580200e-01,-2.472959607839584351e-01,-2.900235056877136230e-01,1.896430850028991699e-01,-1.007863879203796387e-01,-1.251852791756391525e-02,-1.465859562158584595e-01,1.780878156423568726e-01,-3.120823204517364502e-01,1.291723921895027161e-02,2.176860570907592773e-01,-2.588440179824829102e-01,1.567740589380264282e-01,-8.875314891338348389e-02,1.431114822626113892e-01,-7.927271723747253418e-02,3.734678030014038086e-01,-1.235934048891067505e-01,-1.878392137587070465e-02,1.252547651529312134e-01,-2.495816200971603394e-01,-3.412008658051490784e-02,-9.424415230751037598e-02,2.403475530445575714e-02,-1.271171420812606812e-01,1.004246026277542114e-01,-6.776615977287292480e-02,2.086576633155345917e-02,1.203806698322296143e-01,3.388096392154693604e-01,-2.551321983337402344e-01,1.107488796114921570e-01,2.068736255168914795e-01,9.182673878967761993e-03,3.419673740863800049e-01,-6.619603931903839111e-02,2.504039108753204346e-01,-3.285310044884681702e-02,5.807919055223464966e-02,1.882372051477432251e-01,-1.957231201231479645e-02,3.756548091769218445e-02,-3.771427646279335022e-02,1.001068949699401855e-01,4.796762168407440186e-01,1.538818329572677612e-02,2.116000354290008545e-01,-9.692787379026412964e-02,-1.353429164737462997e-02,-6.424796581268310547e-02,2.652154862880706787e-01,1.283384710550308228e-01,1.138196885585784912e-01,3.664042651653289795e-01,-1.299448609352111816e-01);
    -- output layer weights
    constant w2r : w2r_array := (3.938828408718109131e-01,1.251144986599683762e-02,3.898026645183563232e-01,5.647344589233398438e-01,-1.945071965456008911e-01,3.871822655200958252e-01,-4.092536568641662598e-01,1.354921311140060425e-01,-3.196228444576263428e-01,4.516425728797912598e-01,-3.315006569027900696e-02,-5.853371024131774902e-01,1.352412998676300049e-01,-7.582541704177856445e-01,3.652849495410919189e-01,-2.855713963508605957e-01,-9.030334651470184326e-03,-1.951401978731155396e-01,-7.097837328910827637e-01,-1.194379702210426331e-01,-3.674463331699371338e-01,1.732934117317199707e-01,-1.317590326070785522e-01,-2.346892654895782471e-01,-1.203067079186439514e-01,-9.377752989530563354e-02,1.792648285627365112e-01,-3.686468303203582764e-01,2.376415878534317017e-01,4.908555448055267334e-01,-3.188556134700775146e-01,-1.289697457104921341e-02,-4.625348746776580811e-02,1.663445979356765747e-01,2.150007933378219604e-01,3.567383885383605957e-01,3.150950968265533447e-01,1.640192568302154541e-01,1.292601376771926880e-01,-3.842716217041015625e-01,-1.317618694156408310e-02,3.187104314565658569e-02,3.182893693447113037e-01,7.524237781763076782e-02,1.252939458936452866e-02,-3.694263994693756104e-01,2.363408356904983521e-01,-1.709862649440765381e-01,1.911868005990982056e-01,-3.602138757705688477e-01,1.919498294591903687e-01,-2.849886715412139893e-01,9.659691900014877319e-02,9.924292564392089844e-02,5.919287726283073425e-02,-2.608172595500946045e-01,-2.284796349704265594e-02,-2.861020863056182861e-01,-3.743594512343406677e-02,5.469623208045959473e-02,-2.042135000228881836e-01,4.732239246368408203e-01,-1.079529598355293274e-01,1.748222708702087402e-01,-9.621575474739074707e-02,4.691704511642456055e-01,-1.486862599849700928e-01,2.153688073158264160e-01,1.935614943504333496e-01,-1.613049209117889404e-01,-2.816147208213806152e-01,-4.316582977771759033e-01,-1.689505875110626221e-01,-3.079160861670970917e-02,-1.720847189426422119e-01,-1.650388389825820923e-01,2.130784653127193451e-02,-3.176961839199066162e-02,-2.464182376861572266e-01,-4.176778197288513184e-01,-2.689951062202453613e-01,-3.471171259880065918e-01,-1.021618768572807312e-01,-9.428812563419342041e-02,1.890997290611267090e-01,-2.248281091451644897e-01,-1.848896890878677368e-01,-2.064242810010910034e-01,-2.132070809602737427e-01,2.191697955131530762e-01,3.044016063213348389e-01,-3.182524740695953369e-01,2.762046158313751221e-01,4.290765225887298584e-01,1.631522327661514282e-01,-2.243597805500030518e-01,3.019409477710723877e-01,4.401337504386901855e-01,3.674279749393463135e-01,4.948847591876983643e-01,7.160940766334533691e-02,-1.459405422210693359e-01,-2.436342090368270874e-02,1.100217700004577637e-01,5.113604068756103516e-01,5.167697668075561523e-01,-3.310942649841308594e-01,3.678354322910308838e-01,2.305372059345245361e-01,6.823146343231201172e-02,2.063331305980682373e-01,3.957879543304443359e-01,-2.030792534351348877e-01,4.878533631563186646e-02,2.898414433002471924e-02,4.536028504371643066e-01,3.017041832208633423e-02,-6.168825551867485046e-02,-2.339589446783065796e-01,8.012423664331436157e-02,-5.061827227473258972e-02,-1.025797650218009949e-01,1.535278111696243286e-01,2.358022890985012054e-02,4.853000640869140625e-01,1.578418761491775513e-01,7.856775820255279541e-02,-7.077399641275405884e-02,-2.643293440341949463e-01,3.615424036979675293e-01,7.637841254472732544e-02,5.091565251350402832e-01,2.960530519485473633e-01,-5.881276726722717285e-01,2.103932015597820282e-02,5.251191258430480957e-01,7.412775754928588867e-01,-3.456234037876129150e-01,-7.009201049804687500e-01,2.386162132024765015e-01,-7.597284018993377686e-02,-1.987469792366027832e-01,1.491029411554336548e-01,2.308726459741592407e-01,-1.227784976363182068e-01,-7.262875139713287354e-02,5.429552495479583740e-02,-2.845211885869503021e-02,3.048769831657409668e-01,-1.078466475009918213e-01,-1.080727949738502502e-02,-4.719364345073699951e-01,-3.824877142906188965e-01,1.368025690317153931e-01,1.291320379823446274e-02,-2.074646800756454468e-01,1.015291661024093628e-01,4.261896908283233643e-01,3.433902859687805176e-01,-6.850740313529968262e-02,7.342565059661865234e-02,-6.089047715067863464e-02,-6.278201937675476074e-02,-1.572302877902984619e-01,8.428414911031723022e-02,-1.822388470172882080e-01,6.420017778873443604e-02,2.016832083463668823e-01,-3.591150790452957153e-02,-3.989574685692787170e-02,1.910647004842758179e-02,-1.633984893560409546e-01,1.824965626001358032e-01,1.164872571825981140e-01,5.091008543968200684e-01,4.661773797124624252e-03,9.583215415477752686e-02,-7.123275101184844971e-02,-5.127247422933578491e-02,1.764860451221466064e-01,-2.296456396579742432e-01,-9.734843671321868896e-02,-2.325540930032730103e-01,3.206244111061096191e-02,-2.879615724086761475e-01,1.516763716936111450e-01,-3.748078346252441406e-01,-7.801108527928590775e-03,-3.058928251266479492e-01,1.044443845748901367e-01,-5.146752670407295227e-02,-8.172429800033569336e-01,6.099583953619003296e-02,4.506639242172241211e-01,1.799093186855316162e-01,-5.468589663505554199e-01,-2.840094268321990967e-01,4.442441761493682861e-01,3.579969406127929688e-01,1.931589283049106598e-02);
    constant w2r_imag : w2r_array := (-4.111054241657257080e-01,-2.262347191572189331e-02,2.923126220703125000e-01,3.872921168804168701e-01,-3.135396540164947510e-01,2.876935899257659912e-01,-2.909692227840423584e-01,2.537174820899963379e-01,3.158258497714996338e-01,3.325569927692413330e-01,1.475239396095275879e-01,-4.867682754993438721e-01,-3.477280959486961365e-02,-9.418677091598510742e-01,-2.176368981599807739e-01,-2.574050724506378174e-01,-8.864592760801315308e-02,2.280832976102828979e-01,-5.490753054618835449e-01,-1.341833174228668213e-01,3.208375573158264160e-01,1.310365200042724609e-01,-2.520922124385833740e-01,-4.349251687526702881e-01,-2.528760135173797607e-01,-1.874508559703826904e-01,2.763457894325256348e-01,-2.341974228620529175e-01,-2.624804377555847168e-01,3.650273382663726807e-01,4.526355862617492676e-01,9.795399755239486694e-02,-2.339636683464050293e-01,-4.590627271682024002e-03,-6.335910409688949585e-02,3.775125741958618164e-01,-2.912740111351013184e-01,-1.168657019734382629e-01,3.075826764106750488e-01,-4.177189171314239502e-01,-1.184341963380575180e-02,-6.650267168879508972e-03,2.139235585927963257e-01,-1.124552041292190552e-01,-1.107677221298217773e-01,-4.799374043941497803e-01,3.577992618083953857e-01,-5.666213855147361755e-02,-1.758107393980026245e-01,-4.818071722984313965e-01,-8.553355932235717773e-02,-1.894828975200653076e-01,-7.929404824972152710e-02,-7.496469467878341675e-02,8.927067369222640991e-02,-2.390295863151550293e-01,-5.828796327114105225e-02,3.229299187660217285e-01,1.253432929515838623e-01,3.315712511539459229e-02,1.815149039030075073e-01,4.418721497058868408e-01,-2.118335515260696411e-01,-9.002574719488620758e-03,-2.212826907634735107e-01,3.562203347682952881e-01,-3.453345224261283875e-02,3.325710296630859375e-01,-1.856512874364852905e-01,-2.717288434505462646e-01,3.878717124462127686e-01,-3.298319876194000244e-01,-3.459276854991912842e-01,-2.069462984800338745e-01,3.087697327136993408e-01,-1.391240209341049194e-01,-8.284201472997665405e-02,6.989356875419616699e-02,-8.428157120943069458e-02,-4.515679478645324707e-01,2.397925108671188354e-01,-3.846180438995361328e-01,-2.146498858928680420e-01,-2.795165181159973145e-01,7.802072912454605103e-02,-3.234052360057830811e-01,-6.536158919334411621e-02,-8.266906440258026123e-02,2.178481221199035645e-01,1.183627769351005554e-01,-2.128703445196151733e-01,-1.887038201093673706e-01,1.090731024742126465e-01,2.577642202377319336e-01,-5.887200310826301575e-02,-1.841980963945388794e-01,2.911675870418548584e-01,-4.075073003768920898e-01,5.172336101531982422e-01,4.865726828575134277e-01,-9.327714890241622925e-02,-1.757683306932449341e-01,-1.263148635625839233e-01,-7.433554530143737793e-02,3.858963847160339355e-01,4.204976260662078857e-01,-2.114093601703643799e-01,4.855974018573760986e-01,-2.160771787166595459e-01,-4.070915654301643372e-02,-9.323719888925552368e-02,4.943226277828216553e-01,-3.727720975875854492e-01,-1.251572072505950928e-01,1.162551864981651306e-01,4.765591919422149658e-01,-1.201536785811185837e-02,9.769820421934127808e-02,-7.408212870359420776e-02,5.360100790858268738e-02,2.887142077088356018e-02,-1.248440518975257874e-01,4.854347929358482361e-02,-1.523924320936203003e-01,3.637462556362152100e-01,6.931943446397781372e-02,1.984360516071319580e-01,4.251972213387489319e-02,2.453758269548416138e-01,2.805857658386230469e-01,2.651006914675235748e-02,6.264327764511108398e-01,1.448348909616470337e-01,-7.889564037322998047e-01,9.083035588264465332e-02,5.527008175849914551e-01,7.200915813446044922e-01,3.738118708133697510e-01,-5.646389126777648926e-01,2.158636152744293213e-01,7.032618671655654907e-02,-2.351310104131698608e-01,5.809127166867256165e-02,5.456563457846641541e-02,-2.478720098733901978e-01,-1.961555629968643188e-01,1.897235661745071411e-01,8.319061994552612305e-02,-2.850458323955535889e-01,-2.006219029426574707e-01,9.960685670375823975e-02,-3.497138917446136475e-01,-5.485971570014953613e-01,-4.400334879755973816e-02,1.368466615676879883e-01,-1.514685153961181641e-01,1.070991382002830505e-01,-3.903732597827911377e-01,5.015693306922912598e-01,-8.323434740304946899e-02,-9.061527252197265625e-02,-9.832330048084259033e-02,-1.653238832950592041e-01,-3.381399810314178467e-01,-3.687161207199096680e-02,-2.914890944957733154e-01,1.812358796596527100e-01,3.209395706653594971e-01,4.106855019927024841e-02,-1.552376747131347656e-01,9.731732308864593506e-02,-5.878516659140586853e-02,8.123107254505157471e-03,-5.661775544285774231e-02,-3.641085326671600342e-01,2.872396633028984070e-02,-9.248157031834125519e-03,1.059504970908164978e-01,1.143734976649284363e-01,1.714445203542709351e-01,2.056039422750473022e-01,-1.348753869533538818e-01,-3.351184725761413574e-01,-1.589474529027938843e-01,-3.944577276706695557e-01,3.220164403319358826e-02,-2.451488375663757324e-01,1.102622151374816895e-01,3.272062838077545166e-01,-1.883585355244576931e-03,1.533588320016860962e-01,-6.729794144630432129e-01,-1.075431928038597107e-01,2.802771627902984619e-01,-5.422575026750564575e-02,-4.875320494174957275e-01,-2.861402630805969238e-01,-4.166848957538604736e-01,5.100852251052856445e-01,1.058178953826427460e-02);

--    -- Parameters for input and output processing
--    -- min inputs
--    constant p11r : p1r_array := (0.0000000000, 0.0000000000, 0.0262446812);
--    -- 2/(max inputs - min inputs)
--    constant p12r : p1r_array := (2.0595344830, 2.0796091213, 2.1096287436);
--    -- 1's array
--    constant p13r : p1r_array := (1.0000000000, 1.0000000000, 1.0000000000);

--    -- 1's array
--    constant p21r : p2r_array := (1.0000000000, 1.0000000000, 1.0000000000);
--    -- (max targets - min targets)/2
--    constant p22r : p2r_array := (0.4855466166, 0.4808595951, 0.4740170530);
--    -- min targets
--    constant p23r : p2r_array := (0.0000000000, 0.0000000000, 0.0262446812);

    constant input_1 : input_array := (8.993841736943629428e+00,-1.361941648962787355e+01,-3.037512432433412002e+01,-2.303795553990304867e+01,-5.585096528925715731e+00,-2.497185881676191599e-01,-5.803029365706400711e+00,-7.341281717898349157e+00,-2.539568788921599207e+00,-4.012569465444343342e-02,-1.801431598861262806e+00,-2.611664359719903405e+00,-1.126493884330429074e+00,-2.493010498049982870e-01,-6.802824982113042651e-01,-1.090028207264267524e+00,-1.264009516058086646e+00,-1.366371863577403589e+00,-1.174427325366926178e+00,-1.188550052514133704e+00,-1.729556027582755728e+00,-1.774132320409140595e+00,-1.047815788831448325e+00,-9.387890090670355514e-01,-1.527054651998815515e+00,-1.141273276591196151e+00,8.184924656149394906e-04,-1.081435775911523400e-01,-1.170026140825875860e+00,-1.145478434556138403e+00,-3.830735287732123240e-01,-5.045785503003366035e-01,-6.758378183830484609e-01,3.264284650128974619e-01,7.553220025979416885e-01,-8.375324280599354410e-01,-2.163206076939683697e+00,-1.267446099032879969e+00,-2.113063886813558445e-01,-8.693617920066452065e-01,-1.380690082837565225e+00,-1.944483870301980666e-01,8.367454123275444022e-01,2.702613773950162113e-01,-3.582385669901165248e-01,1.198693179983115753e-01,6.235432834645031619e-01,5.079846569387792554e-01,5.035663166361246113e-01,6.391297919828364815e-01,3.619989779097043670e-01,1.924269929059914119e-01,6.496794126716156637e-01,8.216180237112404861e-01,7.356664538220969440e-02,-6.364758586776440019e-01,-5.704453215491839257e-01,-1.978078847837549392e-01,2.564066860774877332e-01,8.976925099544401654e-01,9.988071102718096839e-01,2.003163596649678024e-01,-1.524087171977560606e-01,6.918222225230183930e-01,1.091738014311071092e+00,-5.816969296064655737e-02,-1.052781622801739481e+00,-4.018461943508668810e-01,6.197289573415709629e-01,5.637429101556068467e-01,1.364335436486998621e-01,2.630280817282644179e-01,4.957464054985378787e-01,4.071107168210316707e-01,2.338230806613900148e-01,-1.011380782463464634e-01,-6.429530579928757206e-01,-7.257879496727528412e-01,-2.070651478827806313e-01,3.954307490280140058e-02,-8.766612070801549361e-02,2.522116656522993550e-01,7.934428651386549181e-01,6.064511683450901636e-01,3.117935127403235196e-01,8.295284122122096315e-01,1.069412989530974745e+00,1.534196622790810483e-01,-1.765532674811252090e-01,1.143768323101963302e+00,1.857489405603804489e+00,6.027049362121141840e-01,-1.708970130146663102e-01,9.691790171264076381e-01,1.418698631458786830e+00,-2.139467895348328152e-01,-1.091738014311198768e+00,4.179863029616330827e-01,1.764551802149358473e+00,1.329740592583350978e+00,9.823279398148929697e-01,1.583717322475827194e+00,1.442240497711236635e+00,4.434986123713182682e-01,5.132110947646000287e-01,1.588605142388943570e+00,1.811704197625558788e+00,1.219172769717318250e+00,1.215870845921857235e+00,1.685444887247462109e+00,1.790784950608051762e+00,1.728767161971753286e+00,1.679909711986198095e+00,1.382610775111128953e+00,1.300261992183025628e+00,1.578550848299324905e+00,1.091726067887230478e+00,2.425444470197999913e-01,1.298725069257747666e+00,3.310816441849380176e+00,2.689953436956999511e+00,1.250843562018154387e+00,4.467990552078707545e+00,9.339137693109710980e+00,7.076533449952545851e+00,9.504191533572663442e-01,3.958777391646210564e+00,1.337907178462359425e+01);
--    constant input_2 : input_array := (0.6220960832, 0.6153051526, 0.6091724511, 0.6037398225, 0.5990299621, 0.5950486695, 0.5917875527, 0.5892269339, 0.5873387467, 0.5860892574);
--    constant input_3 : input_array := (0.5813745283, 0.5757680838, 0.5691906670, 0.5617692649, 0.5536314800, 0.5449017861, 0.5356986698, 0.5261326530, 0.5163051276, 0.5063078855);

    constant input_1_i : input_array := (-6.186515414429433868e+00,-4.419520450242567122e+00,-7.691236692636247874e+00,-9.151855319249369458e+00,-4.296684295379975538e+00,1.388368604295092679e-01,-1.113719326034487089e+00,-2.935670749413523239e+00,-9.605049195824824082e-01,6.278164710343806520e-01,-1.186987147687491584e+00,-2.369609137063936277e+00,-8.204420484489491905e-01,-4.257102835010668218e-01,-2.479110219201369425e+00,-3.135390710222994759e+00,-1.575934663004114666e+00,-1.338750639746853821e+00,-2.682852635717558609e+00,-2.273386107025209490e+00,-2.574582473446546671e-01,1.103369713163886434e-01,-1.101192311321611772e+00,-1.120740982822827192e+00,6.853066289608400474e-02,3.496924464667087173e-01,-3.905336787999291737e-01,-8.287554821998868171e-01,-7.806285679030231517e-01,-5.811247921773019520e-01,-1.039507138734512282e-01,3.623333048292751712e-01,3.639126714370193305e-01,2.956154541999795882e-01,3.375959910491657112e-01,-1.976565336017426233e-01,-9.644316065196636423e-01,-5.866327705375975476e-01,3.946513913513702843e-01,5.093914236868957168e-02,-1.038545559250012795e+00,-7.151489911535944266e-01,2.099065377583894110e-01,-6.254323951777973623e-01,-2.031583651382566025e+00,-1.185735214428556006e+00,6.536236216095749896e-01,2.185211994769416521e-01,-1.629452557329613471e+00,-1.659313812434109359e+00,-2.306882830975368059e-01,5.060503183697717677e-02,-5.413195142860844911e-01,-1.766157711721523249e-01,3.605148004559637354e-01,-6.523504126686334725e-01,-2.197689153786825500e+00,-2.197665086205065954e+00,-9.089900627192841753e-01,-7.919040567114288276e-03,-9.233851063999209963e-02,-6.970161639621504923e-01,-1.192324175196056490e+00,-1.024919137940090597e+00,-3.639126714370306548e-01,-2.208959887751420492e-01,-9.163518833884827242e-01,-1.460439212536673192e+00,-1.185647297522177457e+00,-5.588065138652107411e-01,-9.956852936893237360e-02,-4.320503164031008758e-02,-6.421886905842979498e-01,-1.289489988058941217e+00,-6.777708013598364722e-01,7.628648543353627742e-01,9.030937577796074311e-01,-3.774518761280130641e-01,-8.193280918492816811e-01,-1.227863894292129388e-01,-3.995912676540153141e-01,-1.495667718270253133e+00,-9.420003802808168958e-01,7.982029784052567800e-01,6.474908998277892902e-01,-1.141135240206517132e+00,-1.232202487214039355e+00,5.583277503173535994e-01,1.193948483327530230e+00,2.522279386345550600e-01,9.830435320892150219e-02,9.000478985942539367e-01,7.389376815592902936e-01,-2.751578820443991713e-01,-4.765549131038055997e-01,9.973850694608010770e-02,3.639126714370135574e-01,3.040389011364439398e-01,1.597629730845779861e-01,-3.768214186272498267e-01,-9.471830970712782349e-01,-8.561935863988687778e-01,-5.805405938297953927e-01,-6.262832218348510782e-01,-2.700622020792931011e-01,3.661615810062526233e-01,-2.516561391230308642e-01,-1.625090082596159391e+00,-1.286012395160899935e+00,2.047024367056620164e-01,-3.348769462398235586e-01,-2.369677924342284747e+00,-2.217624255004610134e+00,-2.677882929958745883e-01,-2.258061971179002869e-01,-1.570745292611179789e+00,-7.727707602644744433e-01,1.243821777686497043e+00,1.078484499019579879e+00,-9.439056102456144792e-02,5.193098116351959614e-01,1.225254854505461788e+00,3.268969934181350512e-01,8.527240326013472149e-01,3.368973734196655911e+00,2.038509099485522391e+00,-4.599111491188557999e+00,-8.640396798782184362e+00);
--    constant input_2_i : input_array := (-0.6220960832, -0.6153051526, -0.6091724511, 0.6037398225, 0.5990299621, 0.5950486695, 0.5917875527, 0.5892269339, 0.5873387467, 0.5860892574);
--    constant input_3_i : input_array := (-0.5813745283, -0.5757680838, -0.5691906670, 0.5617692649, 0.5536314800, 0.5449017861, 0.5356986698, 0.5261326530, 0.5163051276, 0.5063078855);


end package nn_package;