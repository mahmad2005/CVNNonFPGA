library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package tan_parameters is
    type input_array is array(0 to 1000) of real;-- input array
    type output_array is array(0 to 1000) of real;-- output array
    
    constant fpinput : input_array :=(-5242879.999,-5232394.239,-5221908.479,-5211422.719,-5200936.959,-5190451.199,-5179965.439,-5169479.679,-5158993.919,-5148508.159,-5138022.399,-5127536.639,-5117050.879,-5106565.119,-5096079.359,-5085593.599,-5075107.839,-5064622.079,-5054136.319,-5043650.559,-5033164.799,-5022679.039,-5012193.279,-5001707.519,-4991221.759,-4980735.999,-4970250.239,-4959764.479,-4949278.719,-4938792.959,-4928307.199,-4917821.439,-4907335.679,-4896849.919,-4886364.159,-4875878.399,-4865392.639,-4854906.879,-4844421.119,-4833935.359,-4823449.599,-4812963.839,-4802478.079,-4791992.319,-4781506.559,-4771020.799,-4760535.039,-4750049.279,-4739563.519,-4729077.759,-4718591.999,-4708106.239,-4697620.479,-4687134.719,-4676648.959,-4666163.199,-4655677.439,-4645191.679,-4634705.919,-4624220.159,-4613734.399,-4603248.639,-4592762.879,-4582277.119,-4571791.359,-4561305.599,-4550819.839,-4540334.079,-4529848.319,-4519362.559,-4508876.799,-4498391.039,-4487905.279,-4477419.519,-4466933.759,-4456447.999,-4445962.239,-4435476.479,-4424990.719,-4414504.959,-4404019.199,-4393533.439,-4383047.679,-4372561.919,-4362076.159,-4351590.399,-4341104.639,-4330618.879,-4320133.119,-4309647.359,-4299161.599,-4288675.839,-4278190.079,-4267704.319,-4257218.559,-4246732.799,-4236247.039,-4225761.279,-4215275.519,-4204789.759,-4194303.999,-4183818.239,-4173332.479,-4162846.719,-4152360.959,-4141875.199,-4131389.439,-4120903.679,-4110417.919,-4099932.159,-4089446.399,-4078960.639,-4068474.879,-4057989.119,-4047503.359,-4037017.599,-4026531.839,-4016046.079,-4005560.319,-3995074.559,-3984588.799,-3974103.039,-3963617.279,-3953131.519,-3942645.759,-3932159.999,-3921674.239,-3911188.479,-3900702.719,-3890216.959,-3879731.199,-3869245.439,-3858759.679,-3848273.919,-3837788.159,-3827302.399,-3816816.639,-3806330.879,-3795845.119,-3785359.359,-3774873.599,-3764387.839,-3753902.079,-3743416.319,-3732930.559,-3722444.799,-3711959.039,-3701473.279,-3690987.519,-3680501.759,-3670015.999,-3659530.239,-3649044.479,-3638558.719,-3628072.959,-3617587.199,-3607101.439,-3596615.679,-3586129.919,-3575644.159,-3565158.399,-3554672.639,-3544186.879,-3533701.119,-3523215.359,-3512729.599,-3502243.839,-3491758.079,-3481272.319,-3470786.559,-3460300.799,-3449815.039,-3439329.279,-3428843.519,-3418357.759,-3407871.999,-3397386.239,-3386900.479,-3376414.719,-3365928.959,-3355443.199,-3344957.439,-3334471.679,-3323985.919,-3313500.159,-3303014.399,-3292528.639,-3282042.879,-3271557.119,-3261071.359,-3250585.599,-3240099.839,-3229614.079,-3219128.319,-3208642.559,-3198156.799,-3187671.039,-3177185.279,-3166699.519,-3156213.759,-3145727.999,-3135242.239,-3124756.479,-3114270.719,-3103784.959,-3093299.199,-3082813.439,-3072327.679,-3061841.919,-3051356.159,-3040870.399,-3030384.639,-3019898.879,-3009413.119,-2998927.359,-2988441.599,-2977955.839,-2967470.079,-2956984.319,-2946498.559,-2936012.799,-2925527.039,-2915041.279,-2904555.519,-2894069.759,-2883583.999,-2873098.239,-2862612.479,-2852126.719,-2841640.959,-2831155.199,-2820669.439,-2810183.679,-2799697.919,-2789212.159,-2778726.399,-2768240.639,-2757754.879,-2747269.119,-2736783.359,-2726297.599,-2715811.839,-2705326.079,-2694840.319,-2684354.559,-2673868.799,-2663383.039,-2652897.279,-2642411.519,-2631925.759,-2621439.999,-2610954.239,-2600468.479,-2589982.719,-2579496.959,-2569011.199,-2558525.439,-2548039.679,-2537553.919,-2527068.159,-2516582.399,-2506096.639,-2495610.879,-2485125.119,-2474639.359,-2464153.599,-2453667.839,-2443182.079,-2432696.319,-2422210.559,-2411724.799,-2401239.039,-2390753.279,-2380267.519,-2369781.759,-2359295.999,-2348810.239,-2338324.479,-2327838.719,-2317352.959,-2306867.199,-2296381.439,-2285895.679,-2275409.919,-2264924.159,-2254438.399,-2243952.639,-2233466.879,-2222981.119,-2212495.359,-2202009.599,-2191523.839,-2181038.079,-2170552.319,-2160066.559,-2149580.799,-2139095.039,-2128609.279,-2118123.519,-2107637.759,-2097151.999,-2086666.239,-2076180.479,-2065694.719,-2055208.959,-2044723.199,-2034237.439,-2023751.679,-2013265.919,-2002780.159,-1992294.399,-1981808.639,-1971322.879,-1960837.119,-1950351.359,-1939865.599,-1929379.839,-1918894.079,-1908408.319,-1897922.559,-1887436.799,-1876951.039,-1866465.279,-1855979.519,-1845493.759,-1835007.999,-1824522.239,-1814036.479,-1803550.719,-1793064.959,-1782579.199,-1772093.439,-1761607.679,-1751121.919,-1740636.159,-1730150.399,-1719664.639,-1709178.879,-1698693.119,-1688207.359,-1677721.599,-1667235.839,-1656750.079,-1646264.319,-1635778.559,-1625292.799,-1614807.039,-1604321.279,-1593835.519,-1583349.759,-1572863.999,-1562378.239,-1551892.479,-1541406.719,-1530920.959,-1520435.199,-1509949.439,-1499463.679,-1488977.919,-1478492.159,-1468006.399,-1457520.639,-1447034.879,-1436549.119,-1426063.359,-1415577.599,-1405091.839,-1394606.079,-1384120.319,-1373634.559,-1363148.799,-1352663.039,-1342177.279,-1331691.519,-1321205.759,-1310719.999,-1300234.239,-1289748.479,-1279262.719,-1268776.959,-1258291.199,-1247805.439,-1237319.679,-1226833.919,-1216348.159,-1205862.399,-1195376.639,-1184890.879,-1174405.119,-1163919.359,-1153433.599,-1142947.839,-1132462.079,-1121976.319,-1111490.559,-1101004.799,-1090519.039,-1080033.279,-1069547.519,-1059061.759,-1048575.999,-1038090.239,-1027604.479,-1017118.719,-1006632.959,-996147.199,-985661.438999999,-975175.679,-964689.919,-954204.159,-943718.399,-933232.639,-922746.879,-912261.119,-901775.359,-891289.599,-880803.839,-870318.079,-859832.319,-849346.559,-838860.799,-828375.039,-817889.279,-807403.519,-796917.759,-786431.999,-775946.239,-765460.478999999,-754974.719,-744488.959,-734003.199,-723517.438999999,-713031.679,-702545.919,-692060.159,-681574.398999999,-671088.639,-660602.879,-650117.119,-639631.359,-629145.599,-618659.839,-608174.079,-597688.319,-587202.559,-576716.799,-566231.039,-555745.279,-545259.519,-534773.759,-524287.999,-513802.239,-503316.479,-492830.719,-482344.959,-471859.199,-461373.438999999,-450887.679,-440401.919,-429916.159,-419430.398999999,-408944.639,-398458.879,-387973.119,-377487.359,-367001.599,-356515.839,-346030.079,-335544.319,-325058.559,-314572.799,-304087.039,-293601.279,-283115.519,-272629.759,-262143.999,-251658.239,-241172.479,-230686.719,-220200.959,-209715.199,-199229.438999999,-188743.679,-178257.919,-167772.159,-157286.398999999,-146800.639,-136314.879,-125829.119,-115343.359,-104857.599,-94371.8389999998,-83886.0790000001,-73400.3190000003,-62914.5589999996,-52428.7989999998,-41943.039,-31457.2790000003,-20971.5189999996,-10485.7589999998,0.001,10485.7609999998,20971.5209999996,31457.2810000003,41943.041,52428.8009999998,62914.5609999996,73400.3210000003,83886.0810000001,94371.8409999999,104857.601,115343.361,125829.121,136314.881,146800.641,157286.400999999,167772.161,178257.921,188743.681,199229.440999999,209715.201,220200.961,230686.721,241172.481,251658.241,262144.001,272629.761,283115.521,293601.281,304087.041,314572.801,325058.561,335544.321,346030.081,356515.841,367001.601,377487.361,387973.121,398458.881,408944.641,419430.400999999,429916.161,440401.921,450887.681,461373.440999999,471859.201,482344.961,492830.721,503316.481,513802.241,524288.001,534773.761,545259.521,555745.281,566231.041,576716.801,587202.561,597688.321,608174.081,618659.841,629145.601,639631.361,650117.121,660602.881,671088.641,681574.400999999,692060.161,702545.921,713031.681,723517.441,734003.201,744488.961,754974.721,765460.481,775946.241,786432.001,796917.761,807403.521,817889.281,828375.041,838860.801,849346.561,859832.321,870318.081,880803.841,891289.601,901775.361,912261.121,922746.881,933232.641,943718.401,954204.161,964689.921,975175.681,985661.441,996147.201,1006632.961,1017118.721,1027604.481,1038090.241,1048576.001,1059061.761,1069547.521,1080033.281,1090519.041,1101004.801,1111490.561,1121976.321,1132462.081,1142947.841,1153433.601,1163919.361,1174405.121,1184890.881,1195376.641,1205862.401,1216348.161,1226833.921,1237319.681,1247805.441,1258291.201,1268776.961,1279262.721,1289748.481,1300234.241,1310720.001,1321205.761,1331691.521,1342177.281,1352663.041,1363148.801,1373634.561,1384120.321,1394606.081,1405091.841,1415577.601,1426063.361,1436549.121,1447034.881,1457520.641,1468006.401,1478492.161,1488977.921,1499463.681,1509949.441,1520435.201,1530920.961,1541406.721,1551892.481,1562378.241,1572864.001,1583349.761,1593835.521,1604321.281,1614807.041,1625292.801,1635778.561,1646264.321,1656750.081,1667235.841,1677721.601,1688207.361,1698693.121,1709178.881,1719664.641,1730150.401,1740636.161,1751121.921,1761607.681,1772093.441,1782579.201,1793064.961,1803550.721,1814036.481,1824522.241,1835008.001,1845493.761,1855979.521,1866465.281,1876951.041,1887436.801,1897922.561,1908408.321,1918894.081,1929379.841,1939865.601,1950351.361,1960837.121,1971322.881,1981808.641,1992294.401,2002780.161,2013265.921,2023751.681,2034237.441,2044723.201,2055208.961,2065694.721,2076180.481,2086666.241,2097152.001,2107637.761,2118123.521,2128609.281,2139095.041,2149580.801,2160066.561,2170552.321,2181038.081,2191523.841,2202009.601,2212495.361,2222981.121,2233466.881,2243952.641,2254438.401,2264924.161,2275409.921,2285895.681,2296381.441,2306867.201,2317352.961,2327838.721,2338324.481,2348810.241,2359296.001,2369781.761,2380267.521,2390753.281,2401239.041,2411724.801,2422210.561,2432696.321,2443182.081,2453667.841,2464153.601,2474639.361,2485125.121,2495610.881,2506096.641,2516582.401,2527068.161,2537553.921,2548039.681,2558525.441,2569011.201,2579496.961,2589982.721,2600468.481,2610954.241,2621440.001,2631925.761,2642411.521,2652897.281,2663383.041,2673868.801,2684354.561,2694840.321,2705326.081,2715811.841,2726297.601,2736783.361,2747269.121,2757754.881,2768240.641,2778726.401,2789212.161,2799697.921,2810183.681,2820669.441,2831155.201,2841640.961,2852126.721,2862612.481,2873098.241,2883584.001,2894069.761,2904555.521,2915041.281,2925527.041,2936012.801,2946498.561,2956984.321,2967470.081,2977955.841,2988441.601,2998927.361,3009413.121,3019898.881,3030384.641,3040870.401,3051356.161,3061841.921,3072327.681,3082813.441,3093299.201,3103784.961,3114270.721,3124756.481,3135242.241,3145728.001,3156213.761,3166699.521,3177185.281,3187671.041,3198156.801,3208642.561,3219128.321,3229614.081,3240099.841,3250585.601,3261071.361,3271557.121,3282042.881,3292528.641,3303014.401,3313500.161,3323985.921,3334471.681,3344957.441,3355443.201,3365928.961,3376414.721,3386900.481,3397386.241,3407872.001,3418357.761,3428843.521,3439329.281,3449815.041,3460300.801,3470786.561,3481272.321,3491758.081,3502243.841,3512729.601,3523215.361,3533701.121,3544186.881,3554672.641,3565158.401,3575644.161,3586129.921,3596615.681,3607101.441,3617587.201,3628072.961,3638558.721,3649044.481,3659530.241,3670016.001,3680501.761,3690987.521,3701473.281,3711959.041,3722444.801,3732930.561,3743416.321,3753902.081,3764387.841,3774873.601,3785359.361,3795845.121,3806330.881,3816816.641,3827302.401,3837788.161,3848273.921,3858759.681,3869245.441,3879731.201,3890216.961,3900702.721,3911188.481,3921674.241,3932160.001,3942645.761,3953131.521,3963617.281,3974103.041,3984588.801,3995074.561,4005560.321,4016046.081,4026531.841,4037017.601,4047503.361,4057989.121,4068474.881,4078960.641,4089446.401,4099932.161,4110417.921,4120903.681,4131389.441,4141875.201,4152360.961,4162846.721,4173332.481,4183818.241,4194304.001,4204789.761,4215275.521,4225761.281,4236247.041,4246732.801,4257218.561,4267704.321,4278190.081,4288675.841,4299161.601,4309647.361,4320133.121,4330618.881,4341104.641,4351590.401,4362076.161,4372561.921,4383047.681,4393533.441,4404019.201,4414504.961,4424990.721,4435476.481,4445962.241,4456448.001,4466933.761,4477419.521,4487905.281,4498391.041,4508876.801,4519362.561,4529848.321,4540334.081,4550819.841,4561305.601,4571791.361,4582277.121,4592762.881,4603248.641,4613734.401,4624220.161,4634705.921,4645191.681,4655677.441,4666163.201,4676648.961,4687134.721,4697620.481,4708106.241,4718592.001,4729077.761,4739563.521,4750049.281,4760535.041,4771020.801,4781506.561,4791992.321,4802478.081,4812963.841,4823449.601,4833935.361,4844421.121,4854906.881,4865392.641,4875878.401,4886364.161,4896849.921,4907335.681,4917821.441,4928307.201,4938792.961,4949278.721,4959764.481,4970250.241,4980736.001,4991221.761,5001707.521,5012193.281,5022679.041,5033164.801,5043650.561,5054136.321,5064622.081,5075107.841,5085593.601,5096079.361,5106565.121,5117050.881,5127536.641,5138022.401,5148508.161,5158993.921,5169479.681,5179965.441,5190451.201,5200936.961,5211422.721,5221908.481,5232394.241,5242880.001);
    constant fpoutput : output_array :=(-1048480.79276885,-1048478.86956448,-1048476.90751244,-1048474.9058281,-1048472.863711,-1048470.78034449,-1048468.65489545,-1048466.48651393,-1048464.27433282,-1048462.0174675,-1048459.71501548,-1048457.36605605,-1048454.96964992,-1048452.52483882,-1048450.03064513,-1048447.4860715,-1048444.89010044,-1048442.24169391,-1048439.53979291,-1048436.78331706,-1048433.97116418,-1048431.10220981,-1048428.17530681,-1048425.18928486,-1048422.14295003,-1048419.03508428,-1048415.86444497,-1048412.62976438,-1048409.32974919,-1048405.96307997,-1048402.52841066,-1048399.02436803,-1048395.4495511,-1048391.80253065,-1048388.08184856,-1048384.28601732,-1048380.41351936,-1048376.46280649,-1048372.43229927,-1048368.32038637,-1048364.12542394,-1048359.84573494,-1048355.47960849,-1048351.02529917,-1048346.48102633,-1048341.84497339,-1048337.1152871,-1048332.29007678,-1048327.36741364,-1048322.34532993,-1048317.22181818,-1048311.99483043,-1048306.66227738,-1048301.22202756,-1048295.6719065,-1048290.00969582,-1048284.23313242,-1048278.3399075,-1048272.32766567,-1048266.19400402,-1048259.93647117,-1048253.55256626,-1048247.03973798,-1048240.39538353,-1048233.6168476,-1048226.70142134,-1048219.6463412,-1048212.44878791,-1048205.10588532,-1048197.61469926,-1048189.97223636,-1048182.17544288,-1048174.22120348,-1048166.10633997,-1048157.82761008,-1048149.38170612,-1048140.76525369,-1048131.97481036,-1048123.00686426,-1048113.85783267,-1048104.52406067,-1048095.00181961,-1048085.28730564,-1048075.37663824,-1048065.26585863,-1048054.95092821,-1048044.42772696,-1048033.69205181,-1048022.73961493,-1048011.56604206,-1048000.16687078,-1047988.53754869,-1047976.67343167,-1047964.56978195,-1047952.2217663,-1047939.62445408,-1047926.77281527,-1047913.66171851,-1047900.28592901,-1047886.64010652,-1047872.71880319,-1047858.5164614,-1047844.02741157,-1047829.24586991,-1047814.16593609,-1047798.78159097,-1047783.08669415,-1047767.07498155,-1047750.74006295,-1047734.07541943,-1047717.07440082,-1047699.73022301,-1047682.03596532,-1047663.98456774,-1047645.5688281,-1047626.78139929,-1047607.61478627,-1047588.06134317,-1047568.11327024,-1047547.76261076,-1047527.00124789,-1047505.82090147,-1047484.21312477,-1047462.1693011,-1047439.68064046,-1047416.73817602,-1047393.33276061,-1047369.45506312,-1047345.09556476,-1047320.24455539,-1047294.8921296,-1047269.02818288,-1047242.64240759,-1047215.72428891,-1047188.2631007,-1047160.24790129,-1047131.66752913,-1047102.51059845,-1047072.76549473,-1047042.42037019,-1047011.46313906,-1046979.88147289,-1046947.66279567,-1046914.79427892,-1046881.26283661,-1046847.05512007,-1046812.15751273,-1046776.55612479,-1046740.23678774,-1046703.18504887,-1046665.38616556,-1046626.82509952,-1046587.4865109,-1046547.35475232,-1046506.41386272,-1046464.64756112,-1046422.03924027,-1046378.5719602,-1046334.22844153,-1046288.99105882,-1046242.84183361,-1046195.76242751,-1046147.73413496,-1046098.73787603,-1046048.75418896,-1045997.76322259,-1045945.74472866,-1045892.67805395,-1045838.54213224,-1045783.31547618,-1045726.97616892,-1045669.50185565,-1045610.86973493,-1045551.05654988,-1045490.03857918,-1045427.79162792,-1045364.29101823,-1045299.51157982,-1045233.42764019,-1045166.01301484,-1045097.24099711,-1045027.08434797,-1044955.51528551,-1044882.50547431,-1044808.02601453,-1044732.04743087,-1044654.53966128,-1044575.47204543,-1044494.81331301,-1044412.53157179,-1044328.59429546,-1044242.96831122,-1044155.61978713,-1044066.5142193,-1043975.61641871,-1043882.89049791,-1043788.29985737,-1043691.80717166,-1043593.37437528,-1043492.96264833,-1043390.53240182,-1043286.04326275,-1043179.45405894,-1043070.7228035,-1042959.80667911,-1042846.66202193,-1042731.24430524,-1042613.50812283,-1042493.40717198,-1042370.89423623,-1042245.9211678,-1042118.43886966,-1041988.39727729,-1041855.74534017,-1041720.43100283,-1041582.40118564,-1041441.60176524,-1041297.97755455,-1041151.47228256,-1041002.02857362,-1040849.58792642,-1040694.09069264,-1040535.47605513,-1040373.68200581,-1040208.64532306,-1040040.30154883,-1039868.58496531,-1039693.42857113,-1039514.76405725,-1039332.52178239,-1039146.63074799,-1038957.01857283,-1038763.61146715,-1038566.33420636,-1038365.11010429,-1038159.86098598,-1037950.50716006,-1037736.96739062,-1037519.15886863,-1037296.99718287,-1037070.39629042,-1036839.26848663,-1036603.52437462,-1036363.07283427,-1036117.82099071,-1035867.67418232,-1035612.53592824,-1035352.30789527,-1035086.88986438,-1034816.17969661,-1034540.07329843,-1034258.46458665,-1033971.24545268,-1033678.30572635,-1033379.53313912,-1033074.81328676,-1032764.02959144,-1032447.06326334,-1032123.79326163,-1031794.0962549,-1031457.84658101,-1031114.91620643,-1030765.17468495,-1030408.48911579,-1030044.72410124,-1029673.74170358,-1029295.40140158,-1028909.56004626,-1028516.07181619,-1028114.78817214,-1027705.55781122,-1027288.22662034,-1026862.6376292,-1026428.63096262,-1025986.04379237,-1025534.71028837,-1025074.46156933,-1024605.12565292,-1024126.5274052,-1023638.48848971,-1023140.82731586,-1022633.35898684,-1022115.895247,-1021588.24442872,-1021050.21139871,-1020501.59750388,-1019942.20051667,-1019371.81457994,-1018790.23015134,-1018197.23394726,-1017592.60888639,-1016976.13403274,-1016347.58453837,-1015706.73158571,-1015053.34232945,-1014387.17983818,-1013708.00303564,-1013015.56664171,-1012309.62111311,-1011589.91258387,-1010856.18280558,-1010108.16908745,-1009345.60423621,-1008568.21649591,-1007775.72948764,-1006967.86214917,-1006144.32867458,-1005304.838454,-1004449.09601333,-1003576.80095415,-1002687.64789375,-1001781.32640545,-1000857.52095909,-999915.910861986,-998956.170200118,-997977.967779892,-996980.967070338,-995964.826145905,-994929.197629896,-993873.728638613,-992798.060726289,-991701.829830888,-990584.666220847,-989446.194442839,-988286.033270665,-987103.795655332,-985899.088676445,-984671.513494985,-983420.665307585,-982146.133302405,-980847.500616715,-979524.344296299,-978176.235256792,-976802.738247077,-975403.411814851,-973977.808274512,-972525.473677473,-971045.947785055,-969538.764044096,-968003.449565421,-966439.52510532,-964846.505050189,-963223.897404492,-961571.20378221,-959887.919401935,-958173.533085791,-956427.527262351,-954649.377973734,-952838.554887062,-950994.521310482,-949116.734213919,-947204.644254793,-945257.695808871,-943275.327006486,-941256.969774319,-939202.04988297,-937109.987000528,-934980.194752375,-932812.080787444,-930605.046851165,-928358.488865336,-926071.797015153,-923744.355843648,-921375.544353773,-918964.736118383,-916511.299398358,-914014.597269137,-911473.987755893,-908888.823977627,-906258.454300419,-903582.222500109,-900859.467934667,-898089.525726489,-895271.726954913,-892405.398859174,-889489.865052089,-886524.445744699,-883508.457982138,-880441.215890962,-877322.030938206,-874150.212202378,-870925.066656656,-867645.899464499,-864312.014287901,-860922.713608503,-857477.299061772,-853975.071784448,-850415.332775435,-846797.383270337,-843120.525129776,-839384.061241674,-835587.295937615,-831729.535423429,-827810.088224089,-823828.265643036,-819783.382235978,-815674.756299238,-811501.710372679,-807263.571757211,-802959.673046875,-798589.352675472,-794151.955477668,-789646.833264495,-785073.34541313,-780430.859470806,-775718.75177269,-770936.40807351,-766083.2241927,-761158.606672789,-756161.97345073,-751092.754541812,-745950.3927358,-740734.344304851,-735444.079722772,-730079.08439511,-724638.859399535,-719122.922235935,-713530.807585591,-707862.068078768,-702116.275070012,-696293.01942038,-690391.912285813,-684412.5859108,-678354.694426426,-672217.914651886,-666001.946898452,-659706.515774884,-653331.370993188,-646876.288173621,-640341.069647755,-633725.545258407,-627029.573155178,-620253.040584312,-613395.864671543,-606457.993196556,-599439.405357667,-592340.112525283,-585160.158982649,-577899.622652416,-570558.615807479,-563137.285764532,-555635.815558787,-548054.424598239,-540393.369295898,-532652.943678344,-524833.479969012,-516935.349144545,-508958.961462618,-500904.766959595,-492773.255916409,-484564.959291072,-476280.449116233,-467920.338860224,-459485.283750084,-450975.981055042,-442393.170329032,-433737.633610817,-425010.195580362,-416211.723670156,-407343.128130236,-398405.362045734,-389399.421305837,-380326.344523122,-371187.212902331,-361983.150057688,-352715.321778014,-343384.935738933,-333993.2411616,-324541.528417464,-315031.128578698,-305463.412914039,-295839.792329874,-286161.716756568,-276430.674480101,-266648.191419251,-256815.830348632,-246935.19006808,-237007.904518959,-227035.641848114,-217020.10342031,-206963.022780149,-196866.164564543,-186731.323366997,-176560.322555035,-166355.013042254,-156117.272016604,-145849.001626602,-135552.127627306,-125228.597987992,-114880.381463566,-104509.466131857,-94117.857899038,-83707.5789754738,-73280.6663244401,-62839.1700861748,-52385.1519798338,-41920.6836859587,-31447.8452121493,-20968.7232446529,-10485.4094886469,0.001,10485.4114886469,20968.7252446529,31447.8472121493,41920.6856859587,52385.1539798338,62839.1720861748,73280.6683244401,83707.5809754738,94117.859899038,104509.468131857,114880.383463566,125228.599987992,135552.129627306,145849.003626602,156117.274016604,166355.015042254,176560.324555035,186731.325366997,196866.166564543,206963.024780149,217020.10542031,227035.643848114,237007.906518959,246935.19206808,256815.832348632,266648.19341925,276430.676480101,286161.718756568,295839.794329874,305463.414914039,315031.130578698,324541.530417464,333993.2431616,343384.937738933,352715.323778014,361983.152057688,371187.214902331,380326.346523122,389399.423305837,398405.364045734,407343.130130236,416211.725670156,425010.197580362,433737.635610817,442393.172329032,450975.983055042,459485.285750084,467920.340860224,476280.451116233,484564.961291072,492773.257916409,500904.768959595,508958.963462618,516935.351144545,524833.481969012,532652.945678344,540393.371295898,548054.426598239,555635.817558787,563137.287764532,570558.617807479,577899.624652416,585160.160982649,592340.114525283,599439.407357668,606457.995196556,613395.866671543,620253.042584312,627029.575155178,633725.547258407,640341.071647755,646876.290173621,653331.372993188,659706.517774884,666001.948898452,672217.916651886,678354.696426426,684412.5879108,690391.914285813,696293.02142038,702116.277070012,707862.070078768,713530.809585591,719122.924235935,724638.861399535,730079.08639511,735444.081722772,740734.346304851,745950.3947358,751092.756541812,756161.97545073,761158.60867279,766083.2261927,770936.41007351,775718.753772691,780430.861470806,785073.34741313,789646.835264495,794151.957477668,798589.354675472,802959.675046875,807263.573757211,811501.712372679,815674.758299238,819783.384235978,823828.267643037,827810.09022409,831729.537423429,835587.297937615,839384.063241674,843120.527129776,846797.385270337,850415.334775436,853975.073784448,857477.301061772,860922.715608503,864312.016287901,867645.901464499,870925.068656656,874150.214202378,877322.032938206,880441.217890962,883508.459982138,886524.447744699,889489.867052089,892405.400859174,895271.728954913,898089.527726489,900859.469934667,903582.22450011,906258.456300419,908888.825977628,911473.989755894,914014.599269137,916511.301398358,918964.738118383,921375.546353774,923744.357843648,926071.799015153,928358.490865336,930605.048851165,932812.082787444,934980.196752375,937109.989000528,939202.05188297,941256.971774319,943275.329006486,945257.697808871,947204.646254793,949116.736213919,950994.523310482,952838.556887062,954649.379973734,956427.529262351,958173.535085791,959887.921401935,961571.20578221,963223.899404492,964846.507050189,966439.52710532,968003.451565421,969538.766044096,971045.949785055,972525.475677474,973977.810274513,975403.413814851,976802.740247077,978176.237256792,979524.346296299,980847.502616715,982146.135302405,983420.667307585,984671.515494985,985899.090676445,987103.797655332,988286.035270665,989446.19644284,990584.668220847,991701.831830888,992798.062726289,993873.730638613,994929.199629896,995964.828145906,996980.969070338,997977.969779892,998956.172200118,999915.912861986,1000857.52295909,1001781.32840545,1002687.64989375,1003576.80295415,1004449.09801333,1005304.840454,1006144.33067458,1006967.86414917,1007775.73148764,1008568.21849591,1009345.60623621,1010108.17108745,1010856.18480558,1011589.91458387,1012309.62311311,1013015.56864171,1013708.00503564,1014387.18183818,1015053.34432945,1015706.73358571,1016347.58653837,1016976.13603274,1017592.61088639,1018197.23594726,1018790.23215134,1019371.81657994,1019942.20251667,1020501.59950388,1021050.21339871,1021588.24642872,1022115.897247,1022633.36098684,1023140.82931586,1023638.49048971,1024126.5294052,1024605.12765292,1025074.46356933,1025534.71228837,1025986.04579237,1026428.63296262,1026862.6396292,1027288.22862034,1027705.55981122,1028114.79017214,1028516.07381619,1028909.56204626,1029295.40340158,1029673.74370358,1030044.72610124,1030408.49111579,1030765.17668495,1031114.91820643,1031457.84858101,1031794.0982549,1032123.79526163,1032447.06526334,1032764.03159144,1033074.81528676,1033379.53513912,1033678.30772635,1033971.24745268,1034258.46658665,1034540.07529843,1034816.18169661,1035086.89186438,1035352.30989527,1035612.53792824,1035867.67618232,1036117.82299071,1036363.07483427,1036603.52637462,1036839.27048663,1037070.39829042,1037296.99918287,1037519.16086863,1037736.96939062,1037950.50916006,1038159.86298598,1038365.11210429,1038566.33620636,1038763.61346715,1038957.02057283,1039146.63274799,1039332.52378239,1039514.76605725,1039693.43057113,1039868.58696531,1040040.30354883,1040208.64732306,1040373.68400581,1040535.47805513,1040694.09269264,1040849.58992642,1041002.03057362,1041151.47428256,1041297.97955455,1041441.60376524,1041582.40318564,1041720.43300283,1041855.74734017,1041988.39927729,1042118.44086966,1042245.92316781,1042370.89623623,1042493.40917198,1042613.51012283,1042731.24630524,1042846.66402193,1042959.80867911,1043070.7248035,1043179.45605894,1043286.04526275,1043390.53440182,1043492.96464833,1043593.37637528,1043691.80917166,1043788.30185737,1043882.89249791,1043975.61841871,1044066.5162193,1044155.62178713,1044242.97031122,1044328.59629546,1044412.53357179,1044494.81531301,1044575.47404543,1044654.54166128,1044732.04943087,1044808.02801453,1044882.50747431,1044955.51728551,1045027.08634797,1045097.24299711,1045166.01501484,1045233.42964019,1045299.51357982,1045364.29301823,1045427.79362792,1045490.04057918,1045551.05854988,1045610.87173493,1045669.50385565,1045726.97816892,1045783.31747618,1045838.54413224,1045892.68005395,1045945.74672866,1045997.76522259,1046048.75618896,1046098.73987603,1046147.73613496,1046195.76442751,1046242.84383361,1046288.99305882,1046334.23044153,1046378.5739602,1046422.04124027,1046464.64956112,1046506.41586272,1046547.35675232,1046587.4885109,1046626.82709952,1046665.38816556,1046703.18704887,1046740.23878774,1046776.55812479,1046812.15951273,1046847.05712007,1046881.26483661,1046914.79627892,1046947.66479567,1046979.88347289,1047011.46513906,1047042.42237019,1047072.76749473,1047102.51259845,1047131.66952913,1047160.24990129,1047188.2651007,1047215.72628891,1047242.64440759,1047269.03018288,1047294.8941296,1047320.24655539,1047345.09756476,1047369.45706312,1047393.33476061,1047416.74017602,1047439.68264046,1047462.1713011,1047484.21512477,1047505.82290147,1047527.00324789,1047547.76461076,1047568.11527024,1047588.06334317,1047607.61678627,1047626.78339929,1047645.5708281,1047663.98656774,1047682.03796532,1047699.73222301,1047717.07640082,1047734.07741943,1047750.74206295,1047767.07698155,1047783.08869415,1047798.78359097,1047814.16793609,1047829.24786991,1047844.02941157,1047858.5184614,1047872.72080319,1047886.64210652,1047900.28792901,1047913.66371851,1047926.77481527,1047939.62645408,1047952.2237663,1047964.57178195,1047976.67543167,1047988.53954869,1048000.16887078,1048011.56804206,1048022.74161493,1048033.69405181,1048044.42972697,1048054.95292821,1048065.26785863,1048075.37863824,1048085.28930564,1048095.00381961,1048104.52606067,1048113.85983267,1048123.00886426,1048131.97681036,1048140.76725369,1048149.38370612,1048157.82961008,1048166.10833998,1048174.22320348,1048182.17744288,1048189.97423636,1048197.61669926,1048205.10788532,1048212.45078791,1048219.6483412,1048226.70342134,1048233.6188476,1048240.39738353,1048247.04173798,1048253.55456626,1048259.93847117,1048266.19600402,1048272.32966567,1048278.3419075,1048284.23513242,1048290.01169582,1048295.6739065,1048301.22402756,1048306.66427738,1048311.99683043,1048317.22381818,1048322.34732993,1048327.36941364,1048332.29207678,1048337.1172871,1048341.84697339,1048346.48302633,1048351.02729917,1048355.48160849,1048359.84773494,1048364.12742394,1048368.32238637,1048372.43429927,1048376.46480649,1048380.41551936,1048384.28801732,1048388.08384856,1048391.80453065,1048395.4515511,1048399.02636803,1048402.53041066,1048405.96507997,1048409.33174919,1048412.63176438,1048415.86644497,1048419.03708428,1048422.14495003,1048425.19128486,1048428.17730681,1048431.10420981,1048433.97316418,1048436.78531706,1048439.54179291,1048442.24369391,1048444.89210044,1048447.4880715,1048450.03264513,1048452.52683882,1048454.97164992,1048457.36805605,1048459.71701548,1048462.0194675,1048464.27633282,1048466.48851393,1048468.65689545,1048470.78234449,1048472.865711,1048474.9078281,1048476.90951244,1048478.87156448,1048480.79476885);
end package;